// Verilog netlist created by Tang Dynasty v5.6.66958
// Wed Feb 15 13:03:38 2023

`timescale 1ns / 1ps
module mc_wrapper
  (
  clk,
  ddr_app_addr,
  ddr_app_cmd,
  ddr_app_en,
  ddr_app_wdf_data,
  ddr_app_wdf_end,
  ddr_app_wdf_mask,
  ddr_app_wdf_wren,
  dfi_rddata_dbi_w,
  dfi_rddata_valid_w,
  dfi_rddata_w,
  init_calib_complete,
  rst,
  ddr_app_rd_data,
  ddr_app_rd_data_end,
  ddr_app_rd_data_valid,
  ddr_app_rdy,
  ddr_app_wdf_rdy,
  dfi_act_n_p,
  dfi_address_p,
  dfi_bank_p,
  dfi_bg_p,
  dfi_cas_n_p,
  dfi_cke_p,
  dfi_cs_n_p,
  dfi_odt_p,
  dfi_ras_n_p,
  dfi_rddata_en_p,
  dfi_reset_n,
  dfi_we_n_p,
  dfi_wrdata_en_p,
  dfi_wrdata_mask_p,
  dfi_wrdata_p
  );

  input clk;
  input [26:0] ddr_app_addr;
  input [2:0] ddr_app_cmd;
  input ddr_app_en;
  input [255:0] ddr_app_wdf_data;
  input ddr_app_wdf_end;
  input [31:0] ddr_app_wdf_mask;
  input ddr_app_wdf_wren;
  input [31:0] dfi_rddata_dbi_w;
  input [15:0] dfi_rddata_valid_w;
  input [255:0] dfi_rddata_w;
  input init_calib_complete;
  input rst;
  output [255:0] ddr_app_rd_data;
  output ddr_app_rd_data_end;
  output ddr_app_rd_data_valid;
  output ddr_app_rdy;
  output ddr_app_wdf_rdy;
  output [3:0] dfi_act_n_p;
  output [55:0] dfi_address_p;
  output [11:0] dfi_bank_p;
  output [7:0] dfi_bg_p;
  output [3:0] dfi_cas_n_p;
  output [3:0] dfi_cke_p;
  output [3:0] dfi_cs_n_p;
  output [3:0] dfi_odt_p;
  output [3:0] dfi_ras_n_p;
  output [15:0] dfi_rddata_en_p;
  output [3:0] dfi_reset_n;
  output [3:0] dfi_we_n_p;
  output [15:0] dfi_wrdata_en_p;
  output [31:0] dfi_wrdata_mask_p;
  output [255:0] dfi_wrdata_p;

  parameter ADDR_WIDTH = 14;
  parameter APP_ADDR_WIDTH = 27;
  parameter APP_DATA_WIDTH = 256;
  parameter APP_MASK_WIDTH = 32;
  parameter BANK_GROUP_WIDTH = 2;
  parameter BANK_WIDTH = 3;
  parameter CKE_WIDTH = 1;
  parameter CL = 7;
  parameter COL_WIDTH = 10;
  parameter CS_WIDTH = 1;
  parameter CWL = 6;
  parameter DM_WIDTH = 4;
  parameter DQS_WIDTH = 4;
  parameter DQ_WIDTH = 32;
  parameter DRAM_TYPE = "DDR3";
  parameter ODT_WIDTH = 1;
  parameter ROW_WIDTH = 14;
  parameter SIMULATION = "TRUE";
  parameter nCK_PER_CLK = 4;
  // localparam DATA_BUF_ADDR_WIDTH = 5;
  // localparam MEM_ADDR_ORDER = "ROW_COLUMN_BANK";
  wire [55:0] al_4152494a;
  wire [55:0] al_f09d84cf;
  wire [11:0] al_8b678b52;
  wire [11:0] al_80bec816;
  wire [3:0] al_33061d84;
  wire [3:0] al_44c9e0a6;
  wire [3:0] al_55586ac1;
  wire [3:0] al_2cf67988;
  wire [3:0] al_ac432c54;
  wire [3:0] al_e84b9bda;
  wire [3:0] al_e5dbfdac;
  wire [3:0] al_49010dd2;
  wire [3:0] al_3d66861c;
  wire [3:0] al_733ec639;
  wire [3:0] al_b99d9508;
  wire [3:0] al_94b2715c;
  wire [23:0] al_4732ba15;
  wire [2:0] al_b4da789e;
  wire [23:0] al_2a9196a6;
  wire [2:0] al_48eb6d34;
  wire [23:0] al_72785055;
  wire [2:0] al_d9b4cc10;
  wire  al_8f66e49d;
  wire  al_d31b0b8f;
  wire  al_eac4076b;
  wire  al_20ccc531;
  wire  al_cc069a1e;
  wire  al_96b41fb2;
  wire  al_6051bc62;
  wire  al_66f9507b;
  wire  al_83946844;
  wire  al_cff749bd;
  wire  al_4edaac38;
  wire  al_638fd104;
  wire  al_955d2d0b;
  wire  al_e65434a9;
  wire  al_cd1bc23c;
  wire  al_761b87c7;
  wire  al_62f041ec;
  wire  al_8370ebfb;
  wire  al_e5820766;
  wire  al_62b064bd;
  wire  al_b7f132ea;
  wire  al_33827427;
  wire  al_8c295dd7;
  wire  al_fdbc6cb0;
  wire  al_d0d67001;
  wire  al_2f53f65;
  wire  al_505af09f;
  wire  al_a7c3fab2;
  wire  al_b030bf9a;
  wire  al_3e22da4d;
  wire  al_ddf7a9aa;
  wire  al_c2f4eaf6;
  wire  al_12509175;
  wire  al_f4c5dfba;
  wire  al_9e51440f;
  wire  al_f9950e01;
  wire  al_6bbf1231;
  wire  al_2b0ac92a;
  wire  al_78f859ca;
  wire  al_5cfcbe8d;
  wire  al_35f5fbe2;
  wire  al_9cac2c36;
  wire  al_b7e8ef76;
  wire  al_3a6224d6;
  wire  al_3235c6b2;
  wire  al_8d9f1a8e;
  wire  al_d81bfd7d;
  wire  al_f3aabbcb;
  wire [5:0] al_41bdf331 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_9f61035a /* synthesis ram_style="dram" */ ;
  wire [5:0] al_4e28198f /* synthesis ram_style="dram" */ ;
  wire [5:0] al_af419986 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_cf0afe9a /* synthesis ram_style="dram" */ ;
  wire [5:0] al_f594a8d9 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_df5cbc72 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_cdd95abd /* synthesis ram_style="dram" */ ;
  wire [5:0] al_c5d3b031 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_79af3182 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_efab6074 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_9d72d808 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_a6fdde80 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_e6b17901 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_57e2199e /* synthesis ram_style="dram" */ ;
  wire [5:0] al_48ac75ce /* synthesis ram_style="dram" */ ;
  wire [5:0] al_74387eee /* synthesis ram_style="dram" */ ;
  wire [5:0] al_c7b20b0 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_ff281ad1 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_effd30c4 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_adfe279 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_eec6554e /* synthesis ram_style="dram" */ ;
  wire [5:0] al_905e5060 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_c58c2706 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_b1296b3 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_62b22b32 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_f62f60e1 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_7b737f75 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_d7fecbad /* synthesis ram_style="dram" */ ;
  wire [5:0] al_8d302088 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_95e9fdd1 /* synthesis ram_style="dram" */ ;
  wire [5:0] al_84027ae7 /* synthesis ram_style="dram" */ ;
  wire [4:0] al_194afe0a;
  wire [4:0] al_5e1dd175;
  wire [4:0] al_511af127;
  wire [4:0] al_71c87c87;
  wire [255:0] al_1952ddef;
  wire [255:0] al_31a3e7af;
  wire [31:0] al_c0f3a3cd;
  wire [6:0] al_4aabc590;
  wire [39:0] al_af133298;
  wire [127:0] al_880499db;
  wire [127:0] al_32e78cf2;
  wire [127:0] al_70931fdb;
  wire [127:0] al_2982a0b8;
  wire [127:0] al_cde313f8;
  wire [127:0] al_e3f231cd;
  wire [127:0] al_b43737f6;
  wire [127:0] al_a1c5f121;
  wire [7:0] al_cc4d831c;
  wire [31:0] al_8679dfa;
  wire [6:0] al_ea19deeb;
  wire [15:0] al_523e9f7a;
  wire [15:0] al_4340e4e7;
  wire [15:0] al_55ed1bfd;
  wire [15:0] al_8ef9bc8c;
  wire [15:0] al_e1aabbd4;
  wire [15:0] al_b0d99cb1;
  wire [15:0] al_4f2a09ff;
  wire [15:0] al_f949a7ee;
  wire [4:0] al_5d5ab475;
  wire [0:3] al_d549f91e;
  wire [0:3] al_d7619b2;
  wire [4:0] al_47a64ed5;
  wire [4:0] al_75c1ef4c;
  wire [4:0] al_ce7d4278;
  wire [4:0] al_ad4756a7;
  wire [4:0] al_f8f25e7b;
  wire [4:0] al_3ee9f2ae;
  wire [4:0] al_1f23ce73;
  wire [4:0] al_abc55d75;
  wire [4:0] al_1bc63bd7;
  wire [4:0] al_c2a06982;
  wire [4:0] al_c3bcd0f7;
  wire [4:0] al_35348eec;
  wire [4:0] al_cd4b89ad;
  wire [3:0] al_10206333;
  wire [4:0] al_20b2d1cd;
  wire [1:0] al_b37f6146;
  wire [1:0] al_ffbe21a4;
  wire [1:0] al_d5c3e265;
  wire [3:0] al_73f8a8a7;
  wire [3:0] al_845e0bd1;
  wire [1:0] al_765e8240;
  wire [48:0] al_f0482f12;
  wire [48:0] al_4b620bb0;
  wire [48:0] al_a5104c4f;
  wire [48:0] al_dac85437;
  wire [48:0] al_71f78ff1;
  wire [3:0] al_80083fda;
  wire [4:0] al_dd6ebfb0;
  wire [1:0] al_31adf876;
  wire [4:0] al_b6b411a2;
  wire [2:0] al_a67dc86a;
  wire [2:0] al_c4e56ecb;
  wire [2:0] al_f0abb8e8;
  wire [2:0] al_c46598af;
  wire [2:0] al_7c5b4e5e;
  wire [48:0] al_58851aab;
  wire [3:0] al_c2faf058;
  wire [3:0] al_b5844352;
  wire [3:0] al_a65f5154;
  wire [3:0] al_56b3021d;
  wire [3:0] al_cf91271d;
  wire [4:0] al_81f91ff1;
  wire [4:0] al_7711fc3;
  wire [5:0] al_4213cfc;
  wire [48:0] al_77634075;
  wire [48:0] al_b9ba8b6c;
  wire [48:0] al_9c434c4a;
  wire [48:0] al_d3350acc;
  wire [1:0] al_a9ec6721;
  wire [3:0] al_5453b759;
  wire [48:0] al_b93da8d5;
  wire [48:0] al_6be20a95;
  wire [1:0] al_99c445b5;
  wire [1:0] al_879aba03;
  wire [1:0] al_e484293d;
  wire [48:0] al_3e489598;
  wire [4:0] al_cf086b44;
  wire [0:3] al_886f442e;
  wire [0:3] al_dff56698;
  wire [4:0] al_3b57d409;
  wire [4:0] al_fc7c448b;
  wire [4:0] al_d206e68;
  wire [4:0] al_ce0a0d6b;
  wire [4:0] al_526d80ee;
  wire [4:0] al_c58f63f9;
  wire [4:0] al_44b93047;
  wire [4:0] al_4f585ca5;
  wire [4:0] al_b6ac4cff;
  wire [4:0] al_e42ac584;
  wire [4:0] al_96dda245;
  wire [4:0] al_535746d5;
  wire [4:0] al_c8aa6814;
  wire [3:0] al_9119fd7;
  wire [4:0] al_b90e2b30;
  wire [1:0] al_89251c12;
  wire [1:0] al_40b9c486;
  wire [1:0] al_14c34e2f;
  wire [3:0] al_7a6f3e1;
  wire [3:0] al_c8d0e932;
  wire [1:0] al_bfcf9d28;
  wire [48:0] al_8664dd36;
  wire [48:0] al_393e4b3;
  wire [48:0] al_c6ae1e35;
  wire [48:0] al_b56343fc;
  wire [48:0] al_41f34c81;
  wire [3:0] al_79fcd485;
  wire [4:0] al_31a603ae;
  wire [1:0] al_fd46e088;
  wire [4:0] al_8023991e;
  wire [2:0] al_c289c50a;
  wire [2:0] al_57cd6e45;
  wire [2:0] al_4a605a24;
  wire [2:0] al_90c83bf9;
  wire [3:0] al_8a6bb27f;
  wire [3:0] al_a119035a;
  wire [3:0] al_640bf3cc;
  wire [3:0] al_c3cc6453;
  wire [3:0] al_259bb519;
  wire [4:0] al_8278c32;
  wire [4:0] al_afe3d62c;
  wire [5:0] al_637e5e2a;
  wire [48:0] al_1f1a358;
  wire [48:0] al_9840f3f;
  wire [48:0] al_7dc43980;
  wire [48:0] al_198cecf1;
  wire [3:0] al_f21eb389;
  wire [48:0] al_16a767cd;
  wire [48:0] al_17da2162;
  wire [48:0] al_8ed48b41;
  wire [48:0] al_d9af4975;
  wire [1:0] al_bd042336;
  wire [1:0] al_66e5f5b5;
  wire [1:0] al_3612f044;
  wire [4:0] al_21bd4e5d;
  wire [0:3] al_4bc24ece;
  wire [0:3] al_61614b33;
  wire [4:0] al_c0079c57;
  wire [4:0] al_e2c05b54;
  wire [4:0] al_a2f64ded;
  wire [4:0] al_b1db173b;
  wire [4:0] al_ff390a8f;
  wire [4:0] al_fcd9679a;
  wire [4:0] al_7a57f678;
  wire [4:0] al_402dba27;
  wire [4:0] al_73725553;
  wire [4:0] al_ac18355b;
  wire [4:0] al_d0a384c4;
  wire [4:0] al_1e043bfe;
  wire [4:0] al_b0a8403e;
  wire [3:0] al_a83e1130;
  wire [4:0] al_3e345b21;
  wire [1:0] al_e1208a36;
  wire [1:0] al_11a7c870;
  wire [1:0] al_1f1dc264;
  wire [3:0] al_413c0926;
  wire [3:0] al_6779071c;
  wire [1:0] al_b528368c;
  wire [48:0] al_59b0cd05;
  wire [48:0] al_e9ebbe15;
  wire [48:0] al_c5c971b;
  wire [48:0] al_51cc7f19;
  wire [48:0] al_e6e3a9da;
  wire [3:0] al_cfa51fb3;
  wire [4:0] al_527755ec;
  wire [1:0] al_aaf3456;
  wire [4:0] al_46448d9c;
  wire [2:0] al_369e229d;
  wire [2:0] al_edda145c;
  wire [2:0] al_16929b7c;
  wire [2:0] al_1f97cafb;
  wire [2:0] al_9adc03c8;
  wire [3:0] al_86261d41;
  wire [3:0] al_6824a1b1;
  wire [3:0] al_6d285e98;
  wire [3:0] al_579d2a90;
  wire [3:0] al_2f1f444b;
  wire [4:0] al_7fb24d41;
  wire [4:0] al_e048ecc8;
  wire [5:0] al_e3f59f84;
  wire [48:0] al_31adc4ab;
  wire [48:0] al_39d4ac28;
  wire [48:0] al_2697e1b1;
  wire [48:0] al_f0541159;
  wire [3:0] al_ef92c438;
  wire [48:0] al_8c934a6b;
  wire [48:0] al_4084a330;
  wire [48:0] al_8941a5fb;
  wire [48:0] al_bc0d6480;
  wire [1:0] al_864a13d9;
  wire [1:0] al_f2dedfad;
  wire [1:0] al_ca7553ae;
  wire [4:0] al_f6114766;
  wire [0:3] al_71faa803;
  wire [0:3] al_9c4fa309;
  wire [4:0] al_89ad3a7d;
  wire [4:0] al_45d9e18e;
  wire [4:0] al_c5e4c82d;
  wire [4:0] al_9892447e;
  wire [4:0] al_2497ff95;
  wire [4:0] al_b671fee2;
  wire [4:0] al_c325b022;
  wire [4:0] al_6f7a76fc;
  wire [4:0] al_1a25e1aa;
  wire [4:0] al_dd768853;
  wire [4:0] al_eec54698;
  wire [4:0] al_ffdc699f;
  wire [4:0] al_f1974c03;
  wire [3:0] al_69c2ff54;
  wire [4:0] al_a3f7dedc;
  wire [1:0] al_eacb80c;
  wire [1:0] al_a196b5f4;
  wire [1:0] al_68f1a7a7;
  wire [3:0] al_b25d0e99;
  wire [3:0] al_696c7934;
  wire [1:0] al_e11b20ed;
  wire [48:0] al_974136cc;
  wire [48:0] al_fea7bbd9;
  wire [48:0] al_16b7523e;
  wire [48:0] al_f82ace94;
  wire [48:0] al_7040e81f;
  wire [3:0] al_9941ff24;
  wire [4:0] al_553ae5af;
  wire [1:0] al_4ed70d21;
  wire [4:0] al_5b784e0e;
  wire [2:0] al_9d2be50d;
  wire [2:0] al_7db277fb;
  wire [2:0] al_10aff3dd;
  wire [2:0] al_4795b95a;
  wire  al_cc5fd2c8;
  wire [3:0] al_251b6a5;
  wire [3:0] al_a8314aee;
  wire [3:0] al_ff167b71;
  wire [3:0] al_74d1b04e;
  wire [3:0] al_9d7bf9ff;
  wire [4:0] al_7054a209;
  wire [4:0] al_ba0505cb;
  wire [5:0] al_e6d81dbe;
  wire [48:0] al_3c07b31a;
  wire [48:0] al_fbcce8b0;
  wire [48:0] al_2422b44d;
  wire [48:0] al_9c80d3c6;
  wire [3:0] al_f001c0eb;
  wire [48:0] al_d6e945fd;
  wire [48:0] al_f152e67e;
  wire [48:0] al_ef35f7b6;
  wire [48:0] al_786f2a14;
  wire [1:0] al_b1a73cf;
  wire [1:0] al_1124d2df;
  wire [1:0] al_a1373d93;
  wire [39:0] al_2602b5cf;
  wire [7:0] al_d76fa964;
  wire [3:0] al_90d84dc7;
  wire [3:0] al_a8be2de9;
  wire [1:0] al_a91e0413;
  wire [4:0] al_ee18df00;
  wire [4:0] al_71a56a93;
  wire [4:0] al_f05e4262;
  wire [3:0] al_c360bf4c;
  wire  al_f436c091;
  wire  al_72131b80;
  wire  al_becbe1a2;
  wire  al_4c923ed;
  wire  al_43250e7c;
  wire  al_adcb2e1b;
  wire  al_a2d1acac;
  wire  al_ab3d1147;
  wire  al_d4979c57;
  wire [1:0] al_bc9b7e1e;
  wire [1:0] al_aa505777;
  wire [1:0] al_984f095b;
  wire [1:0] al_1692563a;
  wire [1:0] al_d53ceeb6;
  wire [3:0] al_7ead2bfc;
  wire [7:0] al_53bb123b;
  wire [7:0] al_cbeafa67;
  wire [1:0] al_ef3696df;
  wire  al_b14bdbb3;
  wire  al_9fccc935;
  wire  al_b905b88f;
  wire  al_ccd9a7ea;
  wire  al_e7ffa4ec;
  wire  al_f01dcc55;
  wire  al_ab817290;
  wire [3:0] al_187c11ca;
  wire  al_ac2fd07f;
  wire [1:0] al_437ca69f;
  wire [3:0] al_90a0fe97;
  wire  al_a4894768;
  wire  al_6a408c69;
  wire  al_b8b95ad1;
  wire [3:0] al_81cbac46;
  wire [3:0] al_81c227e0;
  wire  al_12e98266;
  wire  al_68fdf79b;
  wire  al_1c8bee0c;
  wire  al_b05701c2;
  wire  al_826c84b0;
  wire  al_f3fd3c4c;
  wire  al_efe155a8;
  wire  al_d3ca11f1;
  wire  al_9b281de6;
  wire  al_9115a3ab;
  wire  al_a2a57eb6;
  wire  al_8fe5c542;
  wire [7:0] al_eb9aa630;
  wire [7:0] al_3c0a4ef0;
  wire [7:0] al_ecc8e317;
  wire [7:0] al_c8b553c9;
  wire [7:0] al_92812db2;
  wire [7:0] al_534b111d;
  wire [7:0] al_39691102;
  wire [7:0] al_304bc4cf;
  wire [7:0] al_421a630e;
  wire [7:0] al_2cee9b7b;
  wire [7:0] al_2f77b9ea;
  wire [7:0] al_b7a66cc8;
  wire [7:0] al_bce3182d;
  wire [7:0] al_636a0d93;
  wire [7:0] al_e3639d7e;
  wire [7:0] al_18fbbb0f;
  wire [7:0] al_779bd70c;
  wire [7:0] al_45d6e796;
  wire [7:0] al_56820b3e;
  wire [143:0] al_95504971;
  wire [23:0] al_dc65c0d1;
  wire [31:0] al_16ace516;
  wire [9:0] al_c37fabd5;
  wire [2:0] al_9ffa2c81;
  wire [2:0] al_5a67a09b;
  wire [1:0] al_147f1ed5;
  wire [1:0] al_ac2c2542;
  wire [3:0] al_2e186afc;
  wire [3:0] al_c3b79934;
  wire [15:0] al_e736aaf7;
  wire [15:0] al_9f02b6ff;
  wire [15:0] al_a25915f6;
  wire [15:0] al_b340bc6d;
  wire [3:0] al_1d853c9a;
  wire [3:0] al_da91be3;
  wire [3:0] al_887856fc;
  wire [3:0] al_d99aae4d;
  wire [3:0] al_a8d985cf;
  wire [3:0] al_f4295ad6;
  wire [8:0] al_5e053069;
  wire [8:0] al_d07272c1;
  wire [8:0] al_582cdf5;
  wire [8:0] al_a3070745;
  wire [8:0] al_6c3719db;
  wire [8:0] al_fd291354;
  wire [8:0] al_7861e435;
  wire [8:0] al_9c26f92c;
  wire [3:0] al_82fe8ddf;
  wire [3:0] al_92b55720;
  wire [3:0] al_93b093ad;
  wire [3:0] al_8d73b4c8;
  wire [8:0] al_52b895b5;
  wire [8:0] al_bd6aead3;
  wire [8:0] al_febad4d6;
  wire [8:0] al_c57192d3;
  wire [8:0] al_dedaebcb;
  wire [8:0] al_6fe26a79;
  wire [8:0] al_910cb5e3;
  wire [8:0] al_7b9547a0;
  wire [3:0] al_e39e8b51;
  wire [3:0] al_6ad27cba;
  wire [3:0] al_efc928b8;
  wire [3:0] al_d0f70b25;
  wire [9:0] al_c58e2364;
  wire [9:0] al_97b2c696;
  wire [0:0] al_d9786abc;
  wire [0:0] al_72e5ab2f;
  wire [0:0] al_79090ab6;
  wire  al_cc80b352;
  wire  al_c7a09c4f;
  wire [3:0] al_2f365000;
  wire [4:0] al_c9543684;
  wire [3:0] al_cf11b78b;
  wire [3:0] al_9941dfb9;
  wire [3:0] al_b4db00cd;
  wire [14:0] al_48a3872d;
  wire [14:0] al_55d92da7;
  wire [15:0] al_a923bd8;
  wire [3:0] al_bc505469;
  wire [3:0] al_df310708;
  wire [3:0] al_a769a364;
  wire [3:0] al_8b4486c6;
  wire [15:0] al_e827ceba;
  wire [16:0] al_4a27c86;
  wire [0:0] al_c5fa5405;
  wire [0:0] al_dcd8888a;
  wire [3:0] al_a26c7aae;
  wire [26:0] al_58fb4752;
  wire [26:0] al_cf00ed6f;
  wire [26:0] al_5d3f410a;
  wire [2:0] al_88a8db2c;
  wire [2:0] al_65621cdc;
  wire [2:0] al_bfd664bf;
  wire [4:0] al_75c0d27f;
  wire [5:0] al_69b84ba6;
  wire [3:0] al_da88ced7 /* synthesis keep=true */ ;
  wire [5:0] al_3ab36424;
  wire [5:0] al_a3fa002d;
  wire [5:0] al_f3aa16a9;
  wire [5:0] al_d0d403d6;
  wire [5:0] al_2c2ca002;
  wire [5:0] al_5c25a985;
  wire [5:0] al_8b88a45c;
  wire [5:0] al_d88fcc0f;
  wire [5:0] al_b8da42f7;
  wire [5:0] al_f033fc44;
  wire [5:0] al_3a9b666;
  wire [5:0] al_a5ad4b3c;
  wire [5:0] al_77d19440;
  wire [5:0] al_b9ca6681;
  wire [5:0] al_69204309;
  wire [5:0] al_98058573;
  wire [5:0] al_63020263;
  wire [5:0] al_b7a189;
  wire [5:0] al_c527aa4e;
  wire [5:0] al_407652d9;
  wire [5:0] al_fce7b5a9;
  wire [5:0] al_87305132;
  wire [5:0] al_ed19afe1;
  wire [5:0] al_98c6a23b;
  wire [5:0] al_33614149;
  wire [5:0] al_175c7e02;
  wire [5:0] al_b48e0e9a;
  wire [5:0] al_92e7eeea;
  wire [5:0] al_a6a612a6;
  wire [5:0] al_9427b946;
  wire [5:0] al_9bc4f0be;
  wire [5:0] al_764d3602;
  wire [5:0] al_5a84549;
  wire [5:0] al_e5342096;
  wire [5:0] al_c0d076bb;
  wire [5:0] al_27ec7185;
  wire [5:0] al_ea67686c;
  wire [5:0] al_b04b1b3b;
  wire [5:0] al_d55b2543;
  wire [5:0] al_5577a41;
  wire [5:0] al_b0408eb;
  wire [5:0] al_6b6ef69;
  wire [5:0] al_4c1bada4;
  wire [42:0] al_326d3b34 /* synthesis keep=true */ ;
  wire [5:0] al_5362aaf;
  wire [5:0] al_b5082a19;
  wire [5:0] al_d6b9e41;
  wire [5:0] al_4206b0c2;
  wire [5:0] al_44864e28;
  wire [5:0] al_71242bdd;
  wire [5:0] al_100c2219;
  wire [5:0] al_2d22d77a;
  wire [5:0] al_8af537d6;
  wire [5:0] al_175608a7;
  wire [5:0] al_f5e6b3f5;
  wire [5:0] al_abd25e4c;
  wire [5:0] al_9cdd3a01;
  wire [5:0] al_55ef04c8;
  wire [5:0] al_384dd51d;
  wire [5:0] al_269b6545;
  wire [5:0] al_430dd919;
  wire [5:0] al_5c6ba19f;
  wire [5:0] al_4f6bae56;
  wire [5:0] al_206e4ef2;
  wire [5:0] al_ead25ba5;
  wire [5:0] al_b04a4cbc;
  wire [5:0] al_6b9e1d84;
  wire [5:0] al_c244bf8b;
  wire [5:0] al_d44a73a0;
  wire [5:0] al_37663fe4;
  wire [5:0] al_e865b87a;
  wire [5:0] al_f359f0c8;
  wire [5:0] al_85a14e36;
  wire [5:0] al_e31889d8;
  wire [5:0] al_8349e0d1;
  wire [5:0] al_2ef171e7;
  wire [5:0] al_662b3089;
  wire [5:0] al_4a30bd0f;
  wire [5:0] al_2119f32d;
  wire [5:0] al_d9591ec3;
  wire [5:0] al_1d102248;
  wire [5:0] al_f78383db;
  wire [5:0] al_d9be1f39;
  wire [5:0] al_1e255230;
  wire [5:0] al_d61bccef;
  wire [5:0] al_46e8788c;
  wire [5:0] al_56e72bf4;
  wire [42:0] al_57f9dbc3 /* synthesis keep=true */ ;
  wire [4:0] al_aa09a9e5;
  wire [4:0] al_4c8ce587;
  wire [4:0] al_3854534a;
  wire [4:0] al_49eb8970;
  wire [4:0] al_39c7f0b5;
  wire [4:0] al_886fd669;
  wire [4:0] al_3550db07;
  wire [4:0] al_9823c42b;
  wire [4:0] al_90b3a908;
  wire [4:0] al_61edc911;
  wire [4:0] al_abb88584;
  wire [4:0] al_3fe9a5bb;
  wire [4:0] al_e94a3a72;
  wire [4:0] al_57782f22;
  wire [4:0] al_9f1bb485;
  wire [4:0] al_52fa7a1e;
  wire [4:0] al_b81cf447;
  wire [4:0] al_5fdc2ca7;
  wire [4:0] al_2ad878de;
  wire [4:0] al_9ef91e29;
  wire [4:0] al_b1ca7bde;
  wire [4:0] al_54ef982d;
  wire [4:0] al_84ba38ec;
  wire [4:0] al_8bf0a0c9;
  wire [4:0] al_cb2afcca;
  wire [4:0] al_43333b4e;
  wire [4:0] al_ad11f805;
  wire [4:0] al_e4f3a09c;
  wire [4:0] al_eb6aa70a;
  wire [4:0] al_6101d7c8;
  wire [4:0] al_9bd5fcab;
  wire [4:0] al_c408b364;
  wire [4:0] al_b96545cc;
  wire [4:0] al_556b029f;
  wire [4:0] al_4f1aa340;
  wire [4:0] al_902090d1;
  wire [4:0] al_2e33811d;
  wire [4:0] al_6ab65bb5;
  wire [4:0] al_8abfbd08;
  wire [4:0] al_1a0d603f;
  wire [4:0] al_8f8431f6;
  wire [4:0] al_91916c28;
  wire [4:0] al_27625f51;
  wire [42:0] al_a0e1d396 /* synthesis keep=true */ ;
  wire [5:0] al_620ff4d8;
  wire [5:0] al_d62bafb2;
  wire [5:0] al_5d7eff71;
  wire [5:0] al_dd20e4f2;
  wire [257:0] al_955db046;
  wire [3:0] al_2d126bfd;
  wire [4:0] al_17e51133;
  wire [1:0] al_b2febcce;
  wire [1:0] al_4caca369;
  wire [1:0] al_b065182c;
  wire [1:0] al_28515a17;
  wire [1:0] al_19e026e1;
  wire [4:0] al_581e4e41;
  wire [4:0] al_8e42692a;
  wire [4:0] al_7c49eb0a;
  wire [1:0] al_3d403a98;
  wire [4:0] al_b16a7f51;
  wire [4:0] al_880139ce;
  wire [4:0] al_4d6d3de1;
  wire [1:0] al_cc43b80;
  wire [4:0] al_f078a0d3;
  wire [4:0] al_8119a127;
  wire [4:0] al_151512a8;
  wire [1:0] al_16418241;
  wire [4:0] al_cc30604e;
  wire [2:0] al_6b28e3d /* synthesis keep=true */ ;
  wire [4:0] al_dfd53060 /* synthesis keep=true */ ;
  wire [4:0] al_fa928a76 /* synthesis keep=true */ ;
  wire [4:0] al_7b7033c7 /* synthesis keep=true */ ;
  wire [4:0] al_167833a3 /* synthesis keep=true */ ;
  wire [4:0] al_c85123b0 /* synthesis keep=true */ ;
  wire [4:0] al_2b539460 /* synthesis keep=true */ ;
  wire [4:0] al_d23802b0;
  wire [1:0] al_38d9ed4e /* synthesis keep=true */ ;
  wire [1:0] al_6c3e2294 /* synthesis keep=true */ ;
  wire [1:0] al_61432edc /* synthesis keep=true */ ;
  wire [1:0] al_8f9b22bd /* synthesis keep=true */ ;
  wire [1:0] al_a49512ff /* synthesis keep=true */ ;
  wire [1:0] al_d4e10e0d /* synthesis keep=true */ ;
  wire [1:0] al_1719553b;
  wire [1:0] al_9681ccaa;
  wire [1:0] al_1aa44e47;
  wire [1:0] al_f62892;
  wire [2:0] al_7f5f60b /* synthesis keep=true */ ;
  wire [7:0] al_a51937a3 /* synthesis keep=true */ ;
  wire [7:0] al_50ec922d;
  wire [5:0] al_162fb89b;
  wire [255:0] al_c665bb87;
  wire [255:0] al_8235546f;
  wire [31:0] al_e8087d79;
  wire [31:0] al_eb430c3c;
  wire [3:0] al_cdc129c7;
  wire [15:0] al_7cd9f06;
  wire [1:0] al_1e58d748;
  wire [1:0] al_98ae77f2;
  wire [4:0] al_4e964d68;
  wire [3:0] al_57c38d66;
  wire [4:1] al_9c7fabce;
  wire [4:1] al_e0201a;
  wire [287:0] al_3e0d53ab;
  wire [287:0] al_8c7bed02;
  wire [3:0] al_c394d21b;
  wire [3:0] al_a3f66965;
  wire [3:0] al_a2dfc1ad;
  wire [4:0] al_d1db9874;
  wire [4:0] al_3014f961;
  wire al_25e28b94;
  wire al_3c7d7d5c;
  wire al_9ce674e2;
  wire al_e54832a8;
  wire al_29af3518;
  wire al_5c28ad0a;
  wire al_5c9a1fe7;
  wire al_2e89ec2c;
  wire al_754a5a85;
  wire al_a66b7d92;
  wire al_27347df6;
  wire al_4706c253;
  wire al_865f57bc;
  wire al_d273ec64;
  wire al_99e96d3e;
  wire al_53e4871;
  wire al_fa88c9b1;
  wire al_51a8d212;
  wire al_5c8dc62;
  wire al_317c528a;
  wire al_364a5729;
  wire al_950c19d6;
  wire al_1d5f0c20;
  wire al_e7314734;
  wire al_e0ba4c33;
  wire al_dc901033;
  wire al_1bfd1d5e;
  wire al_c1b01733;
  wire al_8ec42bd1;
  wire al_fd33b43;
  wire al_b5aa848;
  wire al_a1fef711;
  wire al_86e6d7f8;
  wire al_cd4f09bc;
  wire al_80aa352a;
  wire al_86a56c9a;
  wire al_159f33b5;
  wire al_1dd73244;
  wire al_a4f25695;
  wire al_2ccfdf18;
  wire al_e6c456f4;
  wire al_97dc1b67;
  wire al_445ee5b3;
  wire al_44ab4bb8;
  wire al_85b0e5ae;
  wire al_31c39442;
  wire al_c9e6a24c;
  wire al_5b6e3903;
  wire al_1f32b3ce;
  wire al_4a3ec7d2;
  wire al_1867b14e;
  wire al_595cd185;
  wire al_d5c31119;
  wire al_dc426867;
  wire al_21194118;
  wire al_2b6ee4f;
  wire al_fc2a0d6e;
  wire al_74d292d1;
  wire al_7ffa75b1;
  wire al_f76f90ba;
  wire al_3cf942a1;
  wire al_e43903c1;
  wire al_512ab51;
  wire al_f3b1307c;
  wire al_b35f14e0;
  wire al_b4f5cc54;
  wire al_6a36379a;
  wire al_78cdcfba;
  wire al_544aea7e;
  wire al_e9d913;
  wire al_20113785;
  wire al_47c5e497;
  wire al_42911267;
  wire al_8abfdb0b;
  wire al_ce5ae5f4;
  wire al_3190947b;
  wire al_a008bee3;
  wire al_dce011d4;
  wire al_ef04f6d;
  wire al_71c5949d;
  wire al_c721314;
  wire al_b9cde5e3;
  wire al_96bd601f;
  wire al_b1f62da3;
  wire al_42c99835;
  wire al_800799cd;
  wire al_8f1d15d4;
  wire al_c6f34b3;
  wire al_85cc6a5c;
  wire al_2cb11ceb;
  wire al_bea784fd;
  wire al_a6b55c3b;
  wire al_6169b199;
  wire al_d83b8ffa;
  wire al_26eb28a;
  wire al_4ccae77b;
  wire al_f33298c;
  wire al_b178800e;
  wire al_ef27da32;
  wire al_ecb49f56;
  wire al_1eef59d6;
  wire al_40c57b0a;
  wire al_f212ca88;
  wire al_7dedd4af;
  wire al_db2237d8;
  wire al_688f86d6;
  wire al_f9d8d0e0;
  wire al_59351be4;
  wire al_697eb2f9;
  wire al_144891ce;
  wire al_5c66c844;
  wire al_d3983157;
  wire al_52ab1d02;
  wire al_3fceb593;
  wire al_2789af72;
  wire al_c803837c;
  wire al_ba93203f;
  wire al_1aca5917;
  wire al_ca5bdee2;
  wire al_806b722b;
  wire al_d1caf9b1;
  wire al_30f2f697;
  wire al_cf317014;
  wire al_196ba081;
  wire al_ba9d658c;
  wire al_3f65b31b;
  wire al_40a2a02d;
  wire al_db637163;
  wire al_eaed5f24;
  wire al_d82546f9;
  wire al_242f965e;
  wire al_d0600950;
  wire al_3ce57cf1;
  wire al_8d9fb1d7;
  wire al_fc29ed6b;
  wire al_61f6a76f;
  wire al_3b96714d;
  wire al_f0955a51;
  wire al_c3cbdf31;
  wire al_4b874e94;
  wire al_421da154;
  wire al_27924928;
  wire al_74987791;
  wire al_855b52a9;
  wire al_52e46bbb;
  wire al_8cc23669;
  wire al_1e4cd67c;
  wire al_d477830d;
  wire al_ff1bd228;
  wire al_353ab8af;
  wire al_33e4a93b;
  wire al_d4d15fe6;
  wire al_7bfa51e5;
  wire al_ebef36bd;
  wire al_f98cca52;
  wire al_a5bb1940;
  wire al_5bf1b92d;
  wire al_14abcb2;
  wire al_47108d32;
  wire al_91f0d008;
  wire al_dc467a61;
  wire al_5bce243b;
  wire al_93118b48;
  wire al_ef0d8a39;
  wire al_776135fb;
  wire al_fb7a2d43;
  wire al_4c1ceb3d;
  wire al_2d7d45f8;
  wire al_61210782;
  wire al_c31bffdd;
  wire al_b265eaef;
  wire al_2cea5c50;
  wire al_6263585f;
  wire al_efa11162;
  wire al_fe8d3a5b;
  wire al_849ce6ee;
  wire al_67f1a13d;
  wire al_ef82c7c1;
  wire al_657419a5;
  wire al_462dcba0;
  wire al_13f4f154;
  wire al_1ec9bae4;
  wire al_b87141aa;
  wire al_7ebd1ee0;
  wire al_d735f43c;
  wire al_d79f3cc5;
  wire al_43d25c67;
  wire al_4b9ffcd1;
  wire al_e690950c;
  wire al_55aa5549;
  wire al_435a6ff0;
  wire al_24aa93c3;
  wire al_4368302f;
  wire al_a9a47c58;
  wire al_bbf70a53;
  wire al_53cc11bb;
  wire al_f7d22b96;
  wire al_b7b6339b;
  wire al_d5903b66;
  wire al_f9d6af3f;
  wire al_5d5a8704;
  wire al_b308bcff;
  wire al_e14ba667;
  wire al_55e91735;
  wire al_5edc286b;
  wire al_24cdfb7e;
  wire al_43e9197c;
  wire al_4966891e;
  wire al_d196f7ed;
  wire al_a1b3ef09;
  wire al_3b949dc9;
  wire al_3996c387;
  wire al_7c792e14;
  wire al_40d3ac10;
  wire al_e2d9e8f4;
  wire al_875e77a3;
  wire al_4afe32e3;
  wire al_e841d4f6;
  wire al_7cd375ed;
  wire al_e2b8e4f5;
  wire al_fcebe00e;
  wire al_dc060d66;
  wire al_37f1795f;
  wire al_6f9e8841;
  wire al_bc31a928;
  wire al_e3e845eb;
  wire al_2be8e99;
  wire al_3e6bc3ac;
  wire al_59b8f11e;
  wire al_ca9ad4fa;
  wire al_7b20e638;
  wire al_b39f3a2d;
  wire al_2f8f631b;
  wire al_21e34e90;
  wire al_7e133bf5;
  wire al_ab7128ba;
  wire al_31b7b66;
  wire al_63dade5d;
  wire al_a9bb616f;
  wire al_5083706f;
  wire al_643bfe7d;
  wire al_f6411514;
  wire al_6f628420;
  wire al_95c3862c;
  wire al_4b08729d;
  wire al_153a7598;
  wire al_838dffd7;
  wire al_19acd84f;
  wire al_e097b175;
  wire al_83bf73ec;
  wire al_342187f3;
  wire al_4cf135b8;
  wire al_9aab1a4f;
  wire al_a87038a;
  wire al_37d972e0;
  wire al_b8516693;
  wire al_ef1fe31d;
  wire al_8abdf99c;
  wire al_34945d75;
  wire al_10c16c;
  wire al_d3acc8ad;
  wire al_4030306c;
  wire al_f6ab792b;
  wire al_2192db1e;
  wire al_1551352;
  wire al_64c4b1ee;
  wire al_cf8fae09;
  wire al_6ddecd31;
  wire al_5949896a;
  wire al_ebc69845;
  wire al_698080d7;
  wire al_a8c83515;
  wire al_b7c175ec;
  wire al_a73e260c;
  wire al_12e89d71;
  wire al_d84d421;
  wire al_e1e4e320;
  wire al_fa0877ed;
  wire al_369dae91;
  wire al_dd59d44c;
  wire al_70d8d4e8;
  wire al_f6c5d1c0;
  wire al_54c46837;
  wire al_f679ae98;
  wire al_f486e5f;
  wire al_29e00248;
  wire al_19d71bde;
  wire al_202cea3f;
  wire al_4124b4b4;
  wire al_75463750;
  wire al_97ed8d08;
  wire al_373390f0;
  wire al_e56639b1;
  wire al_786e90e;
  wire al_84d9df21;
  wire al_5c5f6698;
  wire al_23bdcd5d;
  wire al_867a962f;
  wire al_bb6e492e;
  wire al_9bc80d94;
  wire al_f3f27b05;
  wire al_20384508;
  wire al_b25b5a5a;
  wire al_be7ae2e2;
  wire al_cd1b2b40;
  wire al_961ce596;
  wire al_f748f766;
  wire al_76d4d32b;
  wire al_88804612;
  wire al_1975efd7;
  wire al_f59dd527;
  wire al_dc53c2f4;
  wire al_548ecc42;
  wire al_acf97feb;
  wire al_fe36a6e2;
  wire al_a3a81a88;
  wire al_fad9ab0e;
  wire al_4463b457;
  wire al_42b48cc4;
  wire al_aa2163c2;
  wire al_ce58a1e1;
  wire al_2244f12b;
  wire al_5acc3a2f;
  wire al_8d596be2;
  wire al_d31ef303;
  wire al_8b27a255;
  wire al_4a2d2508;
  wire al_790ebcd;
  wire al_4d6aba82;
  wire al_56881e67;
  wire al_1fba6212;
  wire al_70c902df;
  wire al_72d2fdcd;
  wire al_45a1a0f8;
  wire al_f759090a;
  wire al_45d223ab;
  wire al_f9840a37;
  wire al_9841dcd3;
  wire al_d1b0929d;
  wire al_4779567c;
  wire al_c6c76177;
  wire al_95b46020;
  wire al_95467c49;
  wire al_7a04bdba;
  wire al_e3d7dc13;
  wire al_24ea9f76;
  wire al_48c4d402;
  wire al_4d9c76b0;
  wire al_1f7c5f81;
  wire al_8e0772e5 /* synthesis keep=true */ ;
  wire al_4b38e0f3;
  wire al_9120ce24;
  wire al_7d5b642b;
  wire al_98c339b0;
  wire al_8ee904a8;
  wire al_62952198;
  wire al_92e98f85;
  wire al_1e500c02;
  wire al_718bc19f;
  wire al_cfaa4b74;
  wire al_1c7e0f23;
  wire al_80cba1f;
  wire al_2f87218f;
  wire al_2d60bf7c;
  wire al_2b3c55e4;
  wire al_1fe24196;
  wire al_4c2bab56;
  wire al_b325b551;
  wire al_2761bf91;
  wire al_a5d3389d;
  wire al_840aa4cd;
  wire al_6e2c4231;
  wire al_af3006e2;
  wire al_6cdb74d6;
  wire al_6ab92c75;
  wire al_287c07f8;
  wire al_f9b2e036;
  wire al_5341a91c;
  wire al_591ab1d4;
  wire al_b23d9425;
  wire al_a02f02e8;
  wire al_280c0ef0;
  wire al_d2824414;
  wire al_7cad9721;
  wire al_681e3ff2;
  wire al_9fcbbf12;
  wire al_a4d81981;
  wire al_d3154fbb;
  wire al_97784c51;
  wire al_18326672;
  wire al_688aeb95;
  wire al_8cae5877;
  wire al_e769a1ac;
  wire al_a4dd8227;
  wire al_da2e6045;
  wire al_ac3b1637;
  wire al_533b1c82;
  wire al_41ef913c;
  wire al_17bf017e;
  wire al_c952c11c;
  wire al_ac45c87a;
  wire al_83d9c8d2;
  wire al_227f8a62;
  wire al_4d37ff05;
  wire al_5ec2c98e;
  wire al_bbfb7745;
  wire al_f71dba21;
  wire al_267ffb9b;
  wire al_97814ee2;
  wire al_2b60c4d7;
  wire al_f9500eb2;
  wire al_85770a25;
  wire al_457533f2;
  wire al_5f86f74e;
  wire al_e5cd290d;
  wire al_2f21552f;
  wire al_232e33c9;
  wire al_c8afcceb;
  wire al_50f5aee2;
  wire al_370aa1bb;
  wire al_1b8721f8;
  wire al_1f70c9fe;
  wire al_9e92954d;
  wire al_736e37f2;
  wire al_4f668848;
  wire al_9cb32c9b;
  wire al_899fc7f2;
  wire al_e9f106ba;
  wire al_fd00fe9e;
  wire al_1f4c68e6;
  wire al_d17a0773;
  wire al_95538c25;
  wire al_e0aa83ea;
  wire al_c5c92715;
  wire al_72b4a28e;
  wire al_b741880;
  wire al_d177c6b8;
  wire al_bf6feeb3;
  wire al_f31ca00d;
  wire al_37cdc8a1;
  wire al_8ff2e306;
  wire al_993b1b0f;
  wire al_bc420de3;
  wire al_ece57492;
  wire al_3c73e97d;
  wire al_3b11a186;
  wire al_b0e11bf3;
  wire al_9f6af9ba;
  wire al_c7421999;
  wire al_f9833848;
  wire al_4d38737b;
  wire al_640fb7ec;
  wire al_a315f23;
  wire al_25aa754;
  wire al_53b2015;
  wire al_f11e0936;
  wire al_d017e8b1;
  wire al_667181b3 /* synthesis keep=true */ ;
  wire al_a3c26eaf;
  wire al_3ee0d55a;
  wire al_d53d23aa;
  wire al_1f5636ed;
  wire al_22cfe3fb;
  wire al_ba9c6360;
  wire al_7f9b11b5;
  wire al_bdd2644;
  wire al_67a5cae3;
  wire al_e4ce0401;
  wire al_45e379c7;
  wire al_cd1bbfcd;
  wire al_d4376192;
  wire al_b909a17b;
  wire al_fc597f88;
  wire al_518dbdc;
  wire al_a6b3d6e8;
  wire al_8abd3059;
  wire al_9b9e072a;
  wire al_bfc02a10;
  wire al_9f407117;
  wire al_2873e816;
  wire al_d03801fb;
  wire al_634baaae;
  wire al_a96c64c1;
  wire al_fbbc76d0;
  wire al_89c00c3;
  wire al_b4f15053;
  wire al_3f632af4;
  wire al_94133c8a;
  wire al_7546e20f;
  wire al_84824ed8;
  wire al_10737a6f;
  wire al_65b8bca5;
  wire al_c0aba8fb;
  wire al_571561d4;
  wire al_1a076f81;
  wire al_3fbbb328;
  wire al_f9c028af;
  wire al_7bbf72a3;
  wire al_6969681f;
  wire al_f6b9f88c;
  wire al_5f21f5b9;
  wire al_35747c43;
  wire al_d6220c5c;
  wire al_90fdf0b2;
  wire al_e089a5f3;
  wire al_bc77e2de;
  wire al_c9646708;
  wire al_f6d87ba0;
  wire al_9906a30d;
  wire al_2c190380;
  wire al_3629f8f1;
  wire al_a6dad665;
  wire al_374c386b;
  wire al_f15ca799;
  wire al_e990f0b1;
  wire al_49f2a7a7;
  wire al_7f4f4920;
  wire al_b6b5f546;
  wire al_dac0f49d;
  wire al_4f6e0352;
  wire al_445eda9d;
  wire al_96a3d1d4;
  wire al_2770fee0;
  wire al_5d634c36;
  wire al_928fef0c;
  wire al_77bdc2db;
  wire al_38906f51;
  wire al_ad0a7017;
  wire al_95e1b9d1;
  wire al_d66a1017;
  wire al_c304e63a;
  wire al_8ad763a;
  wire al_799f406d;
  wire al_a9c6b32d;
  wire al_445de8c8;
  wire al_748564c9;
  wire al_bb4f41cb;
  wire al_616d30a;
  wire al_e20bf223;
  wire al_70cc7b9e;
  wire al_44b901ea;
  wire al_33769604;
  wire al_3ab8a708;
  wire al_c83b5b3c;
  wire al_3e34cef0;
  wire al_3a2326ef;
  wire al_f27a52ce;
  wire al_b3f14729;
  wire al_c7d73a75;
  wire al_fcdc6bd3;
  wire al_92899c69;
  wire al_3a54c9a1;
  wire al_ac6abfed;
  wire al_10795ff8;
  wire al_c45c98a0;
  wire al_3fe6e16;
  wire al_751ac083;
  wire al_3d802cc7;
  wire al_fd225290;
  wire al_f56597af;
  wire al_cd9ec0c3;
  wire al_538ebf91;
  wire al_2e98876c;
  wire al_4417e3c3;
  wire al_652e3f22;
  wire al_4ba9f27d;
  wire al_693fd6e1;
  wire al_8d59887e;
  wire al_f589c903;
  wire al_1b24326b;
  wire al_8fb41a59;
  wire al_6ce9ade;
  wire al_8afb85c9;
  wire al_8fe2ae6b;
  wire al_1efa2be8;
  wire al_5773cb6a;
  wire al_15ef40b3;
  wire al_63e01e1c;
  wire al_e7da5efa;
  wire al_4cd1569e;
  wire al_77673c37;
  wire al_1affa237;
  wire al_30c9784a;
  wire al_d253498d;
  wire al_3bb37542;
  wire al_bbfc232e;
  wire al_478a8b50;
  wire al_de3eea8a;
  wire al_fbff2df7;
  wire al_6b420938;
  wire al_f2acf56;
  wire al_845e7508;
  wire al_6a20fb79;
  wire al_9fce8b6a;
  wire al_7d8a45fd;
  wire al_40c85aec;
  wire al_28de045;
  wire al_146c01c2;
  wire al_7c3c9bb5;
  wire al_24cee954;
  wire al_2ee87d50;
  wire al_71e16f2b;
  wire al_91632424;
  wire al_59addda8;
  wire al_7a00688b;
  wire al_8a415a42;
  wire al_3b2c2aa;
  wire al_cebaaa2a;
  wire al_891340a1;
  wire al_99c9c113;
  wire al_ac74f6f1;
  wire al_74e913f6;
  wire al_2bb5f88f;
  wire al_ebce8257;
  wire al_45b542b0;
  wire al_81e393a7;
  wire al_fa36ca4c;
  wire al_b79e57b1;
  wire al_49c007fc;
  wire al_1358b03f;
  wire al_648bb7aa;
  wire al_2d3f245b;
  wire al_afe8fb08;
  wire al_5c104e46;
  wire al_ff3a70dc;
  wire al_c56a3e50;
  wire al_4d76e6af;
  wire al_1c1fb07a;
  wire al_c84bba78;
  wire al_d102b3df;
  wire al_d42c904d;
  wire al_7c9229ee;
  wire al_a6e223da;
  wire al_e1f18395;
  wire al_6896ad14;
  wire al_456c110a;
  wire al_b4ecf439;
  wire al_52665bb8;
  wire al_aafc78b6;
  wire al_28a9f919;
  wire al_993745c8;
  wire al_e7604954;
  wire al_c00d3bb;
  wire al_69a88833;
  wire al_9d7e8bc9;
  wire al_e620c305;
  wire al_96a13ff1;
  wire al_edd1cf59;
  wire al_479ec121;
  wire al_df80405c;
  wire al_a4e4c65a;
  wire al_15b16fc6;
  wire al_55b203da;
  wire al_bb796872;
  wire al_56e36fa5;
  wire al_bbcf8fe1;
  wire al_2a1133de;
  wire al_3cb4c24d;
  wire al_3e1f1b94;
  wire al_a3d2c49d;
  wire al_f7bf47b7;
  wire al_27d253fe;
  wire al_57aea336;
  wire al_e51d86f0;
  wire al_7a27ca16;
  wire al_692dd432;
  wire al_dfa7ddb4;
  wire al_4651c92a;
  wire al_504680b8;
  wire al_ebfbad28;
  wire al_98b1e60d;
  wire al_8025a735;
  wire al_b681403c;
  wire al_cc7cc536;
  wire al_e71d5665;
  wire al_93d3d349;
  wire al_e54eae62;
  wire al_b5b02afa;
  wire al_b6d031c2;
  wire al_8bee4cd6;
  wire al_954ec2c7;
  wire al_4969cacc;
  wire al_895da8d;
  wire al_da34749d;
  wire al_1025128c;
  wire al_691a84bb;
  wire al_2d5968ed;
  wire al_8b4f323b;
  wire al_11b8e521;
  wire al_ff98656b;
  wire al_c621ceb7;
  wire al_9cbe46a;
  wire al_9ccb16fd;
  wire al_da6c82d;
  wire al_f68c5dd8;
  wire al_d2b50474;
  wire al_6e677e24;
  wire al_d712b15f;
  wire al_fd39d17d;
  wire al_112c6aa0;
  wire al_acf6f93e;
  wire al_1aabbc67;
  wire al_7f004572;
  wire al_1827053f;
  wire al_2934d890;
  wire al_3d0b7065;
  wire al_176b7b0e;
  wire al_7c2107c8;
  wire al_5f82f20d;
  wire al_dd0180f1;
  wire al_947ff24d;
  wire al_816f1763;
  wire al_d840d9f3;
  wire al_38e5040b;
  wire al_2b09146;
  wire al_eba4eddb;
  wire al_55cda68f;
  wire al_e7ff6740;
  wire al_51ceabf0;
  wire al_3fdd9bd4;
  wire al_724e96cb;
  wire al_f6cbc027;
  wire al_681de671;
  wire al_6d851644;
  wire al_5b2f4c49;
  wire al_ee675012;
  wire al_b56598d;
  wire al_868dabaf;
  wire al_46fc25e7;
  wire al_22d551b1;
  wire al_af3a3adf;
  wire al_80336d41;
  wire al_fe185597;
  wire al_cf63226f;
  wire al_88d2570b;
  wire al_1ea50fd5;
  wire al_cf05798c;
  wire al_627e01b;
  wire al_9a04ce8f;
  wire al_7aadf07;
  wire al_ab1b96f9;
  wire al_122466dd;
  wire al_25fc271e;
  wire al_fb20038d;
  wire al_ffaa6ed4;
  wire al_9384d2a6;
  wire al_5bb79c4f;
  wire al_f0cf2c1b;
  wire al_a0f44394;
  wire al_ae9de7f7;
  wire al_48347124;
  wire al_ddc7a73f;
  wire al_58f4bcca;
  wire al_4c783ffb;
  wire al_b7e2e71f;
  wire al_c34f057a;
  wire al_195fd12;
  wire al_81d476eb;
  wire al_1f586c30;
  wire al_f53cd64f;
  wire al_5c212f53;
  wire al_b6b9db4;
  wire al_b797198c;
  wire al_73f87281;
  wire al_cafe0ec3;
  wire al_67f78c15;
  wire al_a620188b;
  wire al_a5fb3197;
  wire al_38c33a99;
  wire al_5cd3a57d;
  wire al_fccfd8ff;
  wire al_91e55879;
  wire al_699f3bb8;
  wire al_4ce39135;
  wire al_b93ffb04;
  wire al_d8c260df;
  wire al_42cfbe9b;
  wire al_8b71d8b7;
  wire al_79ca7989;
  wire al_3c683e0a;
  wire al_3b14a515;
  wire al_79ced939;
  wire al_865e3224;
  wire al_310a635;
  wire al_b2200d60;
  wire al_be66ece6;
  wire al_1a3d2fd0;
  wire al_f8a12fba;
  wire al_45523d4b;
  wire al_451ab1e2;
  wire al_38fc89af;
  wire al_e5699c1e;
  wire al_e75d1e47;
  wire al_7a20d1b6;
  wire al_2ccb9cac /* synthesis keep=true */ ;
  wire al_18fc9355;
  wire al_86becd21;
  wire al_e69f53ab;
  wire al_5aa41769;
  wire al_83399132;
  wire al_53ec1776;
  wire al_d7c62deb;
  wire al_60f32aa5;
  wire al_be3efaa4;
  wire al_aecd56b;
  wire al_b13009b2;
  wire al_b0d45bcf;
  wire al_1a4dce1b;
  wire al_100e6173;
  wire al_161ea611;
  wire al_cd0e3f19;
  wire al_2e2c5e0e;
  wire al_128dcf82;
  wire al_5b931dce;
  wire al_7393f55f;
  wire al_5ab672a4;
  wire al_8f446276;
  wire al_c7a5b233;
  wire al_79fd4e7c;
  wire al_4f79a2d4;
  wire al_9ea1824f;
  wire al_fd9fbb70;
  wire al_978813a6;
  wire al_bb5bd57a;
  wire al_9e317c87;
  wire al_3799028a;
  wire al_72d179c3;
  wire al_324d8fba;
  wire al_af37d5e4;
  wire al_7ff14cde;
  wire al_9b7ed9ba;
  wire al_12c68610;
  wire al_59d2fcf;
  wire al_ec69184c;
  wire al_bba532bd;
  wire al_709efed6;
  wire al_41779a5c;
  wire al_d6b1e9ef;
  wire al_cff520de;
  wire al_b3e959dd;
  wire al_b7cccbae;
  wire al_db625dc2;
  wire al_f15041ee;
  wire al_5feeb4d9;
  wire al_4b633b4a;
  wire al_ba842b48;
  wire al_aefc71a0;
  wire al_4b666b4a;
  wire al_ac02de78;
  wire al_a89a7f53;
  wire al_d62c6586;
  wire al_c56838c1;
  wire al_5abac53e;
  wire al_6e29173f;
  wire al_ce965e5b;
  wire al_3e8e72a;
  wire al_8c4b2a57;
  wire al_a27e626a;
  wire al_9bbc19f6;
  wire al_709c747d;
  wire al_c7d91c95;
  wire al_ac6ac5f3;
  wire al_553348a;
  wire al_ce2d52c6;
  wire al_c3834b72;
  wire al_4a355d24;
  wire al_12d74399;
  wire al_42951d78;
  wire al_1ca1a962;
  wire al_1cc0dee2;
  wire al_e2e9d990;
  wire al_cabc97d1;
  wire al_42da1f0d;
  wire al_b65fb56b;
  wire al_edb1c8b0;
  wire al_aa1fb1d9;
  wire al_39c11c38;
  wire al_8a6a56f4;
  wire al_48c3548d;
  wire al_e4c850aa;
  wire al_2057cd57;
  wire al_790e0f32;
  wire al_25e1cc7;
  wire al_4db2fe90;
  wire al_c20a9a7e;
  wire al_56be2a2c;
  wire al_58d81d6c;
  wire al_4396fcc1;
  wire al_ef9d2d1b;
  wire al_6237c511;
  wire al_8932a489;
  wire al_d50c8b50;
  wire al_dfc7aeab;
  wire al_ce5f7b78;
  wire al_856e8c85;
  wire al_10f0cebf;
  wire al_4c28a161;
  wire al_7a822c74;
  wire al_ff84082;
  wire al_49045baf;
  wire al_43b9e423;
  wire al_ca5b8a7;
  wire al_69c0e2e6;
  wire al_59c12bba;
  wire al_19756cb7;
  wire al_23659fe5;
  wire al_15aa8dca;
  wire al_891497d5;
  wire al_2182cd10;
  wire al_61973ebe;
  wire al_f8db84b7;
  wire al_786dc891;
  wire al_fbe54a4d;
  wire al_66395a07;
  wire al_a23768c8;
  wire al_be15f9bd;
  wire al_646e2f99;
  wire al_d2a4a6b0;
  wire al_82bab79d;
  wire al_17c7de95;
  wire al_45251641;
  wire al_3b042d56;
  wire al_514e3a7;
  wire al_ef7c15ad;
  wire al_786b0491;
  wire al_5a2ac1a2;
  wire al_d77bb542;
  wire al_9dfaf151;
  wire al_6f281a7f;
  wire al_8d6dd847;
  wire al_d94dff22;
  wire al_f22292ec;
  wire al_ef2f822e;
  wire al_75fd0159;
  wire al_437081f2;
  wire al_f6e750ed;
  wire al_f735a538;
  wire al_bf156068;
  wire al_6158c618;
  wire al_c9ddcee1;
  wire al_cd0bc85d;
  wire al_7b63babf;
  wire al_f66d7bc0;
  wire al_631e0c37;
  wire al_bd4dc0cb;
  wire al_846eafad;
  wire al_3a754a7b;
  wire al_2e8f51d8;
  wire al_e82b7392;
  wire al_7326000a;
  wire al_77041990;
  wire al_1d36bc6d;
  wire al_b0fb8887;
  wire al_a9552c76;
  wire al_4331638;
  wire al_2a6634d6;
  wire al_19e106e3;
  wire al_c54166ab;
  wire al_41e1e6ea;
  wire al_a01620de;
  wire al_27a9ba79;
  wire al_e59c045a;
  wire al_41fff7fc;
  wire al_2acc39d8;
  wire al_27a5f0e3;
  wire al_dc7ca9c3;
  wire al_3b67e711;
  wire al_764705a7;
  wire al_e9b4dc12;
  wire al_fa80f9c4;
  wire al_65940b21;
  wire al_e5dd3f8d;
  wire al_749a40e9;
  wire al_1cf815c1;
  wire al_c74d7793;
  wire al_82bb1e86;
  wire al_3b347f86;
  wire al_c72051a5;
  wire al_1316088;
  wire al_d8e50712;
  wire al_1c962936;
  wire al_833f5c05;
  wire al_e707cc02;
  wire al_464fb058;
  wire al_9d701591;
  wire al_b1edca88;
  wire al_48aee091;
  wire al_3185ed47;
  wire al_2e96480;
  wire al_9264d6ce;
  wire al_e2bcb10;
  wire al_1b6a0af9;
  wire al_5d3dfa86;
  wire al_403fbf52;
  wire al_8287cea7;
  wire al_a4914504;
  wire al_3df83ccd;
  wire al_e2740cd5;
  wire al_fd5ac0c0;
  wire al_bd5f3c97;
  wire al_364b2d93;
  wire al_10d1f7da;
  wire al_bfe0071c;
  wire al_22a3e261;
  wire al_9dee74a8;
  wire al_25de7719;
  wire al_6a2ba50d;
  wire al_55c1f3f8;
  wire al_53439d34;
  wire al_dedd5989;
  wire al_a1d2ac98;
  wire al_61792012;
  wire al_4743871;
  wire al_6bbd7053;
  wire al_e4c2295a;
  wire al_28da8a0d;
  wire al_539c7732;
  wire al_6692b66c;
  wire al_3647cd0;
  wire al_b62c6ace;
  wire al_49d43cfa;
  wire al_c32d8f29;
  wire al_2f5e01b7;
  wire al_2a5fa8c;
  wire al_b4d9e182;
  wire al_34ff0ff5;
  wire al_286587c2;
  wire al_f498aaed;
  wire al_dd9df6a3;
  wire al_26b95353;
  wire al_e1521e17;
  wire al_a448873e;
  wire al_e80539a7;
  wire al_9526df3b;
  wire al_c959a932;
  wire al_fc1936a5;
  wire al_66bed231;
  wire al_a04a63d4;
  wire al_ebe69372;
  wire al_e0a71537;
  wire al_18d4d578;
  wire al_7ab735a9;
  wire al_37a27dff;
  wire al_d1dcebd4;
  wire al_3303cc51;
  wire al_31da793;
  wire al_eae09b27;
  wire al_9bb5b978;
  wire al_70777327;
  wire al_82050a6e /* synthesis keep=true */ ;
  wire al_cbaa3056;
  wire al_eb7b08f0;
  wire al_a2fce1;
  wire al_1d2d788b;
  wire al_f53b3776;
  wire al_c678831f;
  wire al_7f538ee3;
  wire al_55edb257;
  wire al_e355d8ea;
  wire al_1dde650a;
  wire al_254e8e6;
  wire al_cb650584;
  wire al_d87d83a;
  wire al_f16dd8ea;
  wire al_516990df;
  wire al_1af39dee;
  wire al_9d2235cc;
  wire al_81850512;
  wire al_1d4e62f6;
  wire al_221aa358;
  wire al_2dc3e45;
  wire al_86941e27;
  wire al_4eef0b42;
  wire al_6dee9bef;
  wire al_50105215;
  wire al_63714fc7;
  wire al_6d69b644;
  wire al_70c05302;
  wire al_392853fb;
  wire al_ac21ff42;
  wire al_5e53d63d;
  wire al_6e1be86c;
  wire al_3a4ffd2d;
  wire al_2f16accf;
  wire al_1dbbf5ed;
  wire al_69e722f9;
  wire al_7f1ab5ea;
  wire al_e5b96d96;
  wire al_bd7030bd;
  wire al_31640de4;
  wire al_c3c25a23;
  wire al_2aae8bdf;
  wire al_1370261a;
  wire al_5dbbae98;
  wire al_57c1f314;
  wire al_4aab9ab7;
  wire al_2bdc9af8;
  wire al_a6b23c82;
  wire al_51a643c1;
  wire al_b55a64f2;
  wire al_95fc70f6;
  wire al_7103149d;
  wire al_b7ecdcb9;
  wire al_ac0ca30d;
  wire al_cec7db6;
  wire al_374f7117;
  wire al_169c4c39;
  wire al_be7cdff7;
  wire al_50bc751d;
  wire al_37db4e3;
  wire al_4552d084;
  wire al_ea2829c1;
  wire al_e978fc5;
  wire al_a20b0983;
  wire al_467e7732;
  wire al_8b1b352d;
  wire al_7796e47d;
  wire al_a3e40416;
  wire al_8f975858;
  wire al_b47d0925;
  wire al_f4a06276;
  wire al_b7fe498b;
  wire al_d5de0442;
  wire al_9adb60d3;
  wire al_a4dd1877;
  wire al_6f443675;
  wire al_e72ab4a2;
  wire al_90f5a479;
  wire al_6d99a7bb;
  wire al_10853ef5;
  wire al_712e1022;
  wire al_40276cd4;
  wire al_15ca36a;
  wire al_8d431b3f;
  wire al_a0789cd8;
  wire al_94f083a0;
  wire al_630da3b0;
  wire al_9e2903f5;
  wire al_21302b8a;
  wire al_ba1a11d0;
  wire al_79dddfae;
  wire al_c711503f;
  wire al_ca418906;
  wire al_85567015;
  wire al_b3701730;
  wire al_9860067e;
  wire al_ebb9528c;
  wire al_4135f4fc;
  wire al_ddeaf309;
  wire al_165f2734;
  wire al_a70d3eb4;
  wire al_d6f3e78f;
  wire al_a77bd6b4;
  wire al_114b0fe8;
  wire al_7c6fd728;
  wire al_19014a7b;
  wire al_f7f8cb1;
  wire al_32770943;
  wire al_f01cf98;
  wire al_22cea9d;
  wire al_f7e9a10b;
  wire al_1358d298;
  wire al_8e600ada;
  wire al_629fa86a;
  wire al_ad9637b9;
  wire al_3c502065;
  wire al_f419b7f2;
  wire al_55876a5e;
  wire al_9b520651;
  wire al_9c060979;
  wire al_13f9c71c;
  wire al_6ad3f77e;
  wire al_524a1bfd;
  wire al_dfc3cb3c;
  wire al_87136fec;
  wire al_416ad84c;
  wire al_cb0fcfc7;
  wire al_b2365485;
  wire al_7eb31edc;
  wire al_bdded574;
  wire al_8a3c47e1;
  wire al_3a3118b0;
  wire al_d8ecb3f8;
  wire al_d6e5ffe2;
  wire al_c092a1dc;
  wire al_995c4dc4;
  wire al_b7abf9db;
  wire al_7b43c1e;
  wire al_6860fc86;
  wire al_8cddf958;
  wire al_74055ffa;
  wire al_f027c275;
  wire al_cefb896;
  wire al_485702b6;
  wire al_fa2c6203;
  wire al_e6a713a5;
  wire al_2d84af31;
  wire al_a807c60d;
  wire al_3e892816;
  wire al_732fadca;
  wire al_84bf2198;
  wire al_f748e656;
  wire al_5ea47e0d;
  wire al_4ee2ea2f;
  wire al_3f4770be;
  wire al_509bee50;
  wire al_3ec9b0d6;
  wire al_eedba0b4;
  wire al_5a31c994;
  wire al_1a411806;
  wire al_6ea52063;
  wire al_4d29fbf3;
  wire al_f2c5bff2;
  wire al_862761d2;
  wire al_c28589ac;
  wire al_fb5f7a37;
  wire al_cc48041b;
  wire al_cd905f33;
  wire al_3151fa0;
  wire al_a879fe30;
  wire al_bed6ed0d;
  wire al_8fadd979;
  wire al_28335c6e;
  wire al_5134abf1;
  wire al_d7e366bb;
  wire al_e8c2a90e;
  wire al_dd1e54e7;
  wire al_824b4372;
  wire al_748a22bd;
  wire al_6bd11777;
  wire al_19255c36;
  wire al_63204f4;
  wire al_6f5534a0;
  wire al_f1c7f7af;
  wire al_cf38d855;
  wire al_424bd4b9;
  wire al_802e0d75;
  wire al_2010f91b;
  wire al_c906bdb;
  wire al_5c1c29ee;
  wire al_2f7a19ec;
  wire al_41c51f8;
  wire al_b169d8ec;
  wire al_9c4782d2;
  wire al_3d92dfa6;
  wire al_49679814;
  wire al_884f3fa8;
  wire al_13d7dde4;
  wire al_b63d0e11;
  wire al_2819b010;
  wire al_c64ad91c;
  wire al_c81413d1;
  wire al_4aecdf04;
  wire al_2024cd4b;
  wire al_9d99a742;
  wire al_d301de48;
  wire al_ce2e94ee;
  wire al_44e6dfe9;
  wire al_b091346b;
  wire al_e4f5dc3f;
  wire al_c2e0ff4;
  wire al_91bd4a18;
  wire al_4c19e182;
  wire al_46d55200;
  wire al_98c513dd;
  wire al_5ae0756d;
  wire al_5f6a6401;
  wire al_dcf6b718;
  wire al_4e84d779;
  wire al_1001936c;
  wire al_963a39c1;
  wire al_bc5117fe;
  wire al_92d8fd60;
  wire al_126719a0;
  wire al_e8289617;
  wire al_bc7b13ca;
  wire al_1b5b7fb8;
  wire al_316deb29;
  wire al_7e44c8d5;
  wire al_74066232;
  wire al_7eff70ba;
  wire al_9bbade9e;
  wire al_91941257;
  wire al_df5d8efd;
  wire al_c61f1e9a;
  wire al_3f2ddb8a;
  wire al_8fd7f3b8;
  wire al_7059c89d;
  wire al_ed48bce4;
  wire al_6b5d2018;
  wire al_7564e3b0;
  wire al_3f998e21;
  wire al_2115cf8f;
  wire al_f7549f58;
  wire al_f3529ba5;
  wire al_a0f5de0d;
  wire al_3bcdd651;
  wire al_47aa4bf9;
  wire al_5758806f;
  wire al_ffc3eff4;
  wire al_526ace65;
  wire al_3514085d;
  wire al_270372c;
  wire al_56998d64;
  wire al_93070309;
  wire al_965bd4e5;
  wire al_8954e1e7;
  wire al_53334a6 /* synthesis keep=true */ ;
  wire al_4dd68878;
  wire al_5b157bf;
  wire al_8dcb6b40;
  wire al_af2a474d;
  wire al_177ed223;
  wire al_3f896a8c;
  wire al_90420b48;
  wire al_4a34f384;
  wire al_a4747624;
  wire al_60eb3a40;
  wire al_73c5a4c;
  wire al_39f329dd;
  wire al_e76a8396;
  wire al_e5a22863;
  wire al_bf99db4a;
  wire al_e319e994;
  wire al_d244c645;
  wire al_d271b0a3;
  wire al_a59a1785;
  wire al_a639b152;
  wire al_f9cc5188;
  wire al_386e051a;
  wire al_b537e59c;
  wire al_6df2ab59;
  wire al_759a1829;
  wire al_f7a41bbb;
  wire al_a57e41b7;
  wire al_52d7a8c5;
  wire al_61f2ed17;
  wire al_f7d43aab;
  wire al_a7d66e26;
  wire al_fc5dd8f9;
  wire al_eb1ff054;
  wire al_5f8ecffd;
  wire al_bc72c85a;
  wire al_4904896d;
  wire al_3563cff1;
  wire al_465c1e37;
  wire al_e731c778;
  wire al_542b9ee6;
  wire al_2a4334cc;
  wire al_3ef4ff5b;
  wire al_12aaa92f;
  wire al_7b9f0c1d;
  wire al_323b4714;
  wire al_e4d0aba8;
  wire al_8d2646f7;
  wire al_3ebdb95a;
  wire al_22b5c5ea;
  wire al_d70f37f4;
  wire al_2f6c7b59;
  wire al_d7dd86a1;
  wire al_8860002c;
  wire al_5ffe271b;
  wire al_ef43c30e;
  wire al_724c627b;
  wire al_3ea833b1;
  wire al_dafbe78d;
  wire al_398c67e1;
  wire al_a59eb56e;
  wire al_5b4201dc;
  wire al_be2cdb9a;
  wire al_332b9a71;
  wire al_2a694afc;
  wire al_e1f78661;
  wire al_16866029;
  wire al_4577c722;
  wire al_73962c09;
  wire al_87d947b1;
  wire al_5381ba5b;
  wire al_10938478;
  wire al_73e027c6;
  wire al_17aaf618;
  wire al_5d48c7c5;
  wire al_9abe6c71;
  wire al_432fdaf9;
  wire al_d3f078c4;
  wire al_43cdfb95;
  wire al_a96965a6;
  wire al_bb6dcd3;
  wire al_1c4e8451;
  wire al_a3df3136;
  wire al_52be79ea;
  wire al_ea8a5d3e;
  wire al_388ebe26;
  wire al_48b96055;
  wire al_c4726cab;
  wire al_1c8747c7;
  wire al_f4cc2ce5;
  wire al_321810b0;
  wire al_65e4d4e0;
  wire al_465b8d7d;
  wire al_d149d704;
  wire al_21409483;
  wire al_b97c37dd;
  wire al_c088e9dc;
  wire al_82001be8;
  wire al_8e6a6170;
  wire al_fc44176c;
  wire al_3e56391;
  wire al_ec7a421c;
  wire al_dd965664;
  wire al_2af0d594;
  wire al_4c58e022;
  wire al_198de9a1;
  wire al_9a0a15b5;
  wire al_68e89a39;
  wire al_65bd6ac6;
  wire al_7a15bb7a;
  wire al_a26ecd1c;
  wire al_da7de1b7;
  wire al_cce019;
  wire al_31bcb2f7;
  wire al_b887382e;
  wire al_530cb84f;
  wire al_e650be8a;
  wire al_d4f7298c;
  wire al_b1a37b71;
  wire al_12521532;
  wire al_ce2030ae;
  wire al_f5b9a4c5;
  wire al_cb1ca191;
  wire al_4e72a5eb;
  wire al_c307b680;
  wire al_edebd92e;
  wire al_382cf878;
  wire al_dc12b1d7;
  wire al_b59e0dbf;
  wire al_6d82e9d5;
  wire al_a6bfe69c;
  wire al_a09b37ae;
  wire al_6e8781e4;
  wire al_8a0d8763;
  wire al_afc586c3;
  wire al_4c7c6ba3;
  wire al_d1e349fb;
  wire al_5fff4931;
  wire al_ce21c0de;
  wire al_263ba241;
  wire al_50bc0ffd;
  wire al_440bddc2;
  wire al_bbc46aee;
  wire al_932fd4e1;
  wire al_eaa2008b;
  wire al_2112d3be;
  wire al_ceb1b34b;
  wire al_1549e910;
  wire al_d7badb25;
  wire al_c693d245;
  wire al_3bbe144d;
  wire al_3242da44;
  wire al_9c2c924a;
  wire al_ec32a98f;
  wire al_bc6dea5;
  wire al_238af9ad;
  wire al_43f6f764;
  wire al_9609e9f9;
  wire al_c2672a0d;
  wire al_3bdcd136;
  wire al_618346d9;
  wire al_176f9515;
  wire al_1a7e2632;
  wire al_7f2ef1df;
  wire al_a92e1411;
  wire al_d656ab9;
  wire al_43519c87;
  wire al_6748cc6a;
  wire al_1e6583f2;
  wire al_93fe255e;
  wire al_ca609b89;
  wire al_60bb426f;
  wire al_69127009;
  wire al_6a352978;
  wire al_c4e3d21b;
  wire al_666055dd;
  wire al_c30bbc78;
  wire al_d5d22300;
  wire al_b6f81c2e;
  wire al_1e3dbb5f;
  wire al_b4c6b3bd;
  wire al_ef78cbcb;
  wire al_d51c2ed1;
  wire al_1c402ea2;
  wire al_99fcd329;
  wire al_1f4cc6b;
  wire al_1846303e;
  wire al_c20d9298;
  wire al_54588780;
  wire al_a846796e;
  wire al_4a7b60f;
  wire al_86879761;
  wire al_aed918ac;
  wire al_31deb4f1;
  wire al_712d892b;
  wire al_c8887654;
  wire al_48488f01;
  wire al_58ef9f1a;
  wire al_8704f4a0;
  wire al_24e0f545;
  wire al_9d55a7e5;
  wire al_1c83794e;
  wire al_b15eb135;
  wire al_f7077f69;
  wire al_9d5bb698;
  wire al_432e33d4;
  wire al_10ef1903;
  wire al_eaad117a;
  wire al_1abc6e62;
  wire al_c473b6a4;
  wire al_e395c44e;
  wire al_8454367;
  wire al_caa664ee;
  wire al_fd0c8ec3;
  wire al_332c02d0;
  wire al_a8b491ea;
  wire al_781760a2;
  wire al_d17319e5;
  wire al_96a05b;
  wire al_30565995;
  wire al_b71ef602;
  wire al_c0a7db18;
  wire al_89d8cddf;
  wire al_2242adc3;
  wire al_aead4311;
  wire al_beed7bdd;
  wire al_fe8a405;
  wire al_5c032a2f;
  wire al_1a53fdc6;
  wire al_c330002d;
  wire al_c0693577;
  wire al_76e6275e;
  wire al_fb080638;
  wire al_837d8da3;
  wire al_96d05ba4;
  wire al_18e4b32e;
  wire al_12c2377a;
  wire al_ed3799e7;
  wire al_f42e5022;
  wire al_b6bef94;
  wire al_99ca5e59;
  wire al_7af754c1;
  wire al_3a868c71;
  wire al_18e5c731;
  wire al_9650ab3a;
  wire al_a738798f;
  wire al_72b1cb56;
  wire al_b01ab869;
  wire al_a9ad2b6c;
  wire al_a135e827;
  wire al_7fa83c38;
  wire al_c92d59d9;
  wire al_8194720;
  wire al_7a253edf;
  wire al_231ef4df;
  wire al_13a574fa;
  wire al_fb9a605b;
  wire al_db7ff57e;
  wire al_4e6ba179;
  wire al_237c733d;
  wire al_7d5a8c76;
  wire al_9b32a85e;
  wire al_2374b47d;
  wire al_7e2e3620;
  wire al_8dc1b606;
  wire al_35f3cf28;
  wire al_bfe50c52;
  wire al_f149b540;
  wire al_53cd58ac;
  wire al_b3e9d06c;
  wire al_c84ffce0;
  wire al_c5d5a3f6;
  wire al_d46ec896;
  wire al_79f445c4;
  wire al_6b991e1c;
  wire al_5dd540e5;
  wire al_57b41659;
  wire al_2d6bf5be;
  wire al_842732c2;
  wire al_b3d60ef7;
  wire al_fb5f08ff;
  wire al_90254f7;
  wire al_b9ff4892;
  wire al_63860ff5;
  wire al_15578244;
  wire al_21e21c;
  wire al_9602e904;
  wire al_6d6f00e5;
  wire al_c8a2915b;
  wire al_570aaefb;
  wire al_3589ff80;
  wire al_1aea9b48;
  wire al_4483f4ea;
  wire al_9af29299;
  wire al_af82789;
  wire al_37c023d;
  wire al_b5a5e144;
  wire al_9388375e;
  wire al_bf3d0760;
  wire al_8211c6dd;
  wire al_fbec08cf;
  wire al_d3598a31;
  wire al_385080cf;
  wire al_80f00b;
  wire al_484d3915;
  wire al_c9eb9f8c;
  wire al_8c8e8f6a;
  wire al_6f337ab4;
  wire al_2cd04711;
  wire al_f13534df;
  wire al_c48ef761;
  wire al_9e404664;
  wire al_198bf41a;
  wire al_d39ce0c;
  wire al_b71b7f68;
  wire al_4ba8484b;
  wire al_a1fbbbd1;
  wire al_58de2ea4;
  wire al_db15dba5;
  wire al_db39a0bd;
  wire al_c3565be1;
  wire al_6f81b627;
  wire al_76bac341;
  wire al_588f198a;
  wire al_9ac35c50;
  wire al_5606bbf4;
  wire al_c993dae4;
  wire al_a06bb9a1;
  wire al_4b03c837;
  wire al_f8e44d17;
  wire al_ff1cf72f;
  wire al_46b8ac3c;
  wire al_41c9267e;
  wire al_c58b049c;
  wire al_1ffff680;
  wire al_be11f694;
  wire al_f88e71cf;
  wire al_dfdff5e7;
  wire al_a45ee49d;
  wire al_7de91657;
  wire al_2fdead54;
  wire al_73697ad3;
  wire al_482dfbbf;
  wire al_853f0be5;
  wire al_b7fd68ad;
  wire al_d323ca15;
  wire al_7f632198;
  wire al_35c78d09;
  wire al_6e02c90c;
  wire al_6f3fb610;
  wire al_5f022649;
  wire al_21c5d9e6;
  wire al_312cedcc;
  wire al_ba2fb587;
  wire al_f43a0c3c;
  wire al_fd5b02e2;
  wire al_9a41ae4f;
  wire al_b366bb58;
  wire al_6784532f;
  wire al_6c8827e1;
  wire al_8a1c71af;
  wire al_6d9415b;
  wire al_e735abef;
  wire al_2a364bea;
  wire al_1cc7635e;
  wire al_c4e50727;
  wire al_aa8528c4;
  wire al_12af440;
  wire al_174c5495;
  wire al_a6bf875b;
  wire al_1fe9b96a;
  wire al_afe8a6f9;
  wire al_e4885785;
  wire al_1495678c;
  wire al_a807e4d3;
  wire al_66c80cd2;
  wire al_7f9da669;
  wire al_9b835e77;
  wire al_58bba036;
  wire al_90876008;
  wire al_7959b11f;
  wire al_22ec870;
  wire al_484f859d;
  wire al_fc9b7dfa;
  wire al_45d2984c;
  wire al_855245d9;
  wire al_68e325c6;
  wire al_4f00db65;
  wire al_ca978bef;
  wire al_713543ac;
  wire al_c0d8b545;
  wire al_24009166;
  wire al_eec1ba11;
  wire al_dc674b57;
  wire al_6d33eaeb;
  wire al_fa46dbba;
  wire al_a3c61604;
  wire al_7fdd8f7a;
  wire al_b16882ef;
  wire al_20ae9484;
  wire al_3f6a9f97;
  wire al_370abec1;
  wire al_15b509ab;
  wire al_6255d7f7;
  wire al_a082bc48;
  wire al_154c9279;
  wire al_18aca87e;
  wire al_f57af6b4;
  wire al_b2bde781;
  wire al_69c9761a;
  wire al_67ffb718;
  wire al_be5b15b0;
  wire al_685b247;
  wire al_47147006;
  wire al_7b2556ad;
  wire al_698dfed0;
  wire al_1223a962;
  wire al_80311da5;
  wire al_c62e8a82;
  wire al_2d260a04;
  wire al_12563419;
  wire al_e32a2e7c;
  wire al_d31fa142;
  wire al_55232c98;
  wire al_524ab3e2;
  wire al_fbd177b5;
  wire al_bc808160;
  wire al_e29cf77;
  wire al_5ece979a;
  wire al_a76392f;
  wire al_fcb84919;
  wire al_ac3a915e;
  wire al_f100fb27;
  wire al_1f5470a8;
  wire al_b6610a70;
  wire al_5bb559f0;
  wire al_432340bb;
  wire al_3f592f2c;
  wire al_ee2d8b77;
  wire al_54b33a69;
  wire al_2ca74a7;
  wire al_ef9accde;
  wire al_6a03de0;
  wire al_c9d121b2;
  wire al_99917cb7;
  wire al_8514591d;
  wire al_c1a95cc7;
  wire al_4566fdd3;
  wire al_49733697;
  wire al_2957c84b;
  wire al_c79b855c;
  wire al_3ac9505a;
  wire al_ad018368;
  wire al_4bd4fa38;
  wire al_434e6eb1;
  wire al_365f3d23;
  wire al_b0784ca8;
  wire al_badd7923;
  wire al_79c695eb;
  wire al_3a7e0263;
  wire al_9a44af5;
  wire al_4ae2fdc2;
  wire al_3bfb3478;
  wire al_9b29508b;
  wire al_db03633e;
  wire al_fe37e390;
  wire al_743fb5ed;
  wire al_c8295b95;
  wire al_ec4a81f;
  wire al_40d806bd;
  wire al_45a34621;
  wire al_cb5fd325;
  wire al_9680139f;
  wire al_7d50905e;
  wire al_92e38148;
  wire al_eb5035c8;
  wire al_6cc9e68d;
  wire al_ca0e45f8;
  wire al_f44df3e;
  wire al_d7181d37;
  wire al_c3029dcc;
  wire al_3ba0cc79;
  wire al_2d8af247;
  wire al_e3c7998c;
  wire al_eb540174;
  wire al_90b7699;
  wire al_18ebfba6;
  wire al_cb6618b2;
  wire al_8e57b8ea;
  wire al_3225efe4;
  wire al_c18a6fab;
  wire al_a6b572a3;
  wire al_7941134;
  wire al_28570942;
  wire al_4e9593a4;
  wire al_ac57883f;
  wire al_3e848d66;
  wire al_42f2763a;
  wire al_fff872b2;
  wire al_acfaa45c;
  wire al_a83cb045;
  wire al_c1f0ed98;
  wire al_4f7a36e8;
  wire al_c5705f8a;
  wire al_9821c430;
  wire al_898823b1;
  wire al_731b9711;
  wire al_62d3bb1d;
  wire al_21374d40;
  wire al_1cd23aa7;
  wire al_11b28491;
  wire al_aca36a53;
  wire al_813c693b /* synthesis keep=true */ ;
  wire al_7c29888a;
  wire al_4c03fc24;
  wire al_330ee0e3;
  wire al_e58efc01;
  wire al_bf594241;
  wire al_10f4d190;
  wire al_489041e9;
  wire al_61f44420;
  wire al_aab837cc;
  wire al_a7c937ec;
  wire al_66006155;
  wire al_54004a97;
  wire al_5a6db454;
  wire al_1308b999;
  wire al_8dcceed9;
  wire al_adf8e398;
  wire al_355d4013;
  wire al_e4f8f2fd;
  wire al_903070b1;
  wire al_f33f7f41;
  wire al_5ace851;
  wire al_e825eb09;
  wire al_a90a7b11;
  wire al_2ded3658;
  wire al_5068e71b;
  wire al_9ef819de;
  wire al_6b872c5;
  wire al_58e4bd8e;
  wire al_fdaccc20;
  wire al_ce84f7a6;
  wire al_11041b8b;
  wire al_fe081845;
  wire al_9d23d003;
  wire al_a12892b0;
  wire al_ddd2e3de;
  wire al_de2b5681;
  wire al_4830d0fa;
  wire al_b0eff5ca;
  wire al_fd64f6c3;
  wire al_d3947eeb;
  wire al_c6d66579;
  wire al_a9ffc103;
  wire al_7ee48c14;
  wire al_2599c30;
  wire al_1b9ef62a;
  wire al_9ab94adf;
  wire al_799ff6e6;
  wire al_eb0a7105;
  wire al_dd2698f4;
  wire al_793e445;
  wire al_858348d9;
  wire al_e2481062;
  wire al_3f0f44a5;
  wire al_ee9d432a;
  wire al_2eed0a97;
  wire al_264acb9b;
  wire al_ce170fdf;
  wire al_19a0944b;
  wire al_eaa78f2d;
  wire al_7b7614e0;
  wire al_ab431a20;
  wire al_f2d75fa6;
  wire al_ab2d2d18;
  wire al_beea7df8;
  wire al_6694e9cf;
  wire al_a735e2bc;
  wire al_99214f52;
  wire al_5b58c5a7;
  wire al_b578c72c;
  wire al_f0eae58e;
  wire al_ed6ca683;
  wire al_366699aa;
  wire al_cffc4db7;
  wire al_7ee9bd9c;
  wire al_7b5e551b;
  wire al_3613b64a;
  wire al_1c42289;
  wire al_41ff936b;
  wire al_97559555;
  wire al_613310ab;
  wire al_821df217;
  wire al_754cb61b;
  wire al_8f668693;
  wire al_815d1ad6;
  wire al_757240b3;
  wire al_2d8e01f3;
  wire al_8825809e;
  wire al_90caa0c7;
  wire al_1dd9faa9;
  wire al_ce8339bf;
  wire al_18a07add;
  wire al_c3339143;
  wire al_e7e914bb;
  wire al_32c129b3;
  wire al_f5ca45d2;
  wire al_60141953;
  wire al_cf94ebc3;
  wire al_4053f9a0;
  wire al_36161b0f;
  wire al_2775bd20;
  wire al_290f1dfa;
  wire al_57d1b933;
  wire al_45e32f1a;
  wire al_f3161340;
  wire al_2570708b;
  wire al_6f3de2dc;
  wire al_60fd4192;
  wire al_f2987856;
  wire al_ba1ded0d;
  wire al_32460991;
  wire al_a92f34f8;
  wire al_6c74032f;
  wire al_a91a268;
  wire al_14184769;
  wire al_c9258181;
  wire al_478aa8b9;
  wire al_94a7a40;
  wire al_2a63dd17;
  wire al_4704250e;
  wire al_432975cc;
  wire al_dfa5ff6c;
  wire al_d211a035;
  wire al_dc492d87;
  wire al_c37042bd;
  wire al_944bd830;
  wire al_3624cfe0;
  wire al_12dd86af;
  wire al_189dc8c0;
  wire al_9609a6f5;
  wire al_bf0c650;
  wire al_34c94edb;
  wire al_4ca26c83;
  wire al_1a3a4ed7;
  wire al_f60ec0d5;
  wire al_df5418e9;
  wire al_83ae9a40;
  wire al_56102450;
  wire al_ddf07c29;
  wire al_f7a09f99;
  wire al_116d91a8;
  wire al_3197cad9;
  wire al_8f13de6b;
  wire al_dc9abd46;
  wire al_8f5d07af;
  wire al_2a43f573;
  wire al_9752d581;
  wire al_a7c305cd;
  wire al_32307526;
  wire al_ddc0b8a6;
  wire al_ab813978;
  wire al_52694b4b;
  wire al_bd85c50d;
  wire al_13f5c59d;
  wire al_7329b916;
  wire al_21a638b3;
  wire al_3d90e9a3;
  wire al_e377f7a4;
  wire al_7cf355db;
  wire al_b6ed5e1b;
  wire al_63293fc5;
  wire al_5477c30f;
  wire al_aff4e477;
  wire al_e7777d0d;
  wire al_ec64ca16;
  wire al_ebf34b40;
  wire al_aeeedc7e;
  wire al_42eb8568;
  wire al_8ec0a0c8;
  wire al_acd1c245;
  wire al_fd1d15be;
  wire al_7f125c63;
  wire al_61e4c12;
  wire al_e75ba485;
  wire al_594d9eef;
  wire al_f6290e5d;
  wire al_9f34fb19;
  wire al_e96a29f2;
  wire al_e0bee367;
  wire al_ad44d351;
  wire al_27647c5b;
  wire al_359de7f7;
  wire al_84cbc97b;
  wire al_a2e27860;
  wire al_29e29c2;
  wire al_3fb2454f;
  wire al_47d4f942;
  wire al_b7074965;
  wire al_bc75ce6f;
  wire al_4a9b23a9;
  wire al_cee52ae5;
  wire al_ad9326a7;
  wire al_3c305c5d;
  wire al_d77438af;
  wire al_75ba7c3a;
  wire al_cf7de8fd;
  wire al_4cb51ed9;
  wire al_efc69db4;
  wire al_969bce5a;
  wire al_5bb4cdbf;
  wire al_466952a1;
  wire al_6e5cc87d;
  wire al_ce51fefb;
  wire al_875002d2;
  wire al_23ffeaf6;
  wire al_ab1a88b1;
  wire al_b7ba8863;
  wire al_6a0564ce;
  wire al_e8b6474b;
  wire al_f2a9e54d;
  wire al_36fbd71d;
  wire al_800e1ab8;
  wire al_55d82b12;
  wire al_65273b79;
  wire al_199366db;
  wire al_e1e03eb2;
  wire al_7581b68c;
  wire al_e53fc54d;
  wire al_c3b5911e;
  wire al_e9d8781;
  wire al_552a02c8;
  wire al_45ef6b15;
  wire al_322f98e5;
  wire al_2684592f;
  wire al_186881f4;
  wire al_def29dc7;
  wire al_12797435;
  wire al_eb32138;
  wire al_56ab2c31;
  wire al_fdc5c136;
  wire al_f838789f;
  wire al_31c210;
  wire al_36b0c0a;
  wire al_a201d3b2;
  wire al_9a4d5ae0;
  wire al_6bb6f9ee;
  wire al_81f7233;
  wire al_71703480;
  wire al_d7bd990b;
  wire al_739cb624;
  wire al_eeb27c9c;
  wire al_32cf3ccd;
  wire al_bcb724be;
  wire al_581cf91a;
  wire al_ea7f7c64;
  wire al_80d96d10;
  wire al_a98f5d5;
  wire al_696ce813;
  wire al_422c6d68;
  wire al_aec0250a;
  wire al_90969885;
  wire al_5fe1070b;
  wire al_83fb54f8;
  wire al_2039287b;
  wire al_890d7ece;
  wire al_290e28a2;
  wire al_ef0a54ec;
  wire al_a540be99;
  wire al_34ca0b86;
  wire al_70337de1;
  wire al_da48a4d6;
  wire al_d44a1539;
  wire al_5e34a0d9;
  wire al_187efcc;
  wire al_691042b7;
  wire al_eb9d8684;
  wire al_9e7f07bf;
  wire al_6224ca70;
  wire al_77706154;
  wire al_f6e3dfbd;
  wire al_810f7f51;
  wire al_c3077309;
  wire al_ff2cde7a;
  wire al_31adef42;
  wire al_223e27a1;
  wire al_e250e193;
  wire al_c4db602d;
  wire al_177e297a;
  wire al_14d0a20a;
  wire al_a855268a;
  wire al_4476a641;
  wire al_33a1ab04;
  wire al_ebd8858;
  wire al_a0a71833;
  wire al_9cc84a67;
  wire al_80baf9fa;
  wire al_c9b8e286;
  wire al_7038cb56;
  wire al_309702b;
  wire al_401f1215;
  wire al_5d0bc72b;
  wire al_ad7bbe14;
  wire al_bbb63b9;
  wire al_e4a5394c;
  wire al_dac9476c;
  wire al_2f7efa54;
  wire al_85e91cf0;
  wire al_527ad770;
  wire al_50c08ac;
  wire al_163e3e0c;
  wire al_7fda6214;
  wire al_d524c6a5;
  wire al_a6968310;
  wire al_1556ef5b;
  wire al_e0f76854;
  wire al_bbd8d9ee;
  wire al_9f44cd3f;
  wire al_81777b16;
  wire al_f996058d;
  wire al_f1d76027;
  wire al_cdb85e5d;
  wire al_7bd1a9d6;
  wire al_31b57a77;
  wire al_c3f3285c;
  wire al_7d2b45a1;
  wire al_fbacc3a8;
  wire al_b9053852;
  wire al_5fc98ca9;
  wire al_e42e193d;
  wire al_312f6ab1;
  wire al_7b6b3d00;
  wire al_b349d1f9;
  wire al_241ce585;
  wire al_8b91849a;
  wire al_e220508d;
  wire al_ba559767;
  wire al_189beaf8;
  wire al_c4ec8088;
  wire al_7a2b0bb8;
  wire al_ebe8b3b7;
  wire al_920bfd47;
  wire al_fbdfd137;
  wire al_b10901c4;
  wire al_d0e0cc74;
  wire al_7077034d;
  wire al_4d2207ab;
  wire al_b7580b14;
  wire al_84c4e89e;
  wire al_4e77858f;
  wire al_c4cdc14c;
  wire al_c88a646f;
  wire al_a9ba8e79;
  wire al_82ccfd38;
  wire al_956bd9e3;
  wire al_ef3dcd46;
  wire al_74787620;
  wire al_41c60d64;
  wire al_64ae12a2;
  wire al_eaf1b77d;
  wire al_98025056;
  wire al_63db5a9c;
  wire al_785b323e;
  wire al_bfe09e38;
  wire al_46e8cf64;
  wire al_c2d49ea8;
  wire al_ce0ffb93;
  wire al_3c9faf77;
  wire al_a75ec498;
  wire al_3128e6f;
  wire al_9898f5d2;
  wire al_78d64c6e;
  wire al_f06f70db;
  wire al_421f3e11;
  wire al_1df0d799;
  wire al_aa84749f;
  wire al_de545759;
  wire al_2534fd55;
  wire al_3f8224e9;
  wire al_cc0caf5a;
  wire al_748cb5ab;
  wire al_b9ce4338;
  wire al_997d115c;
  wire al_881110e;
  wire al_df8baf16;
  wire al_9cb4bf74;
  wire al_16e3e4ef;
  wire al_320b8e92;
  wire al_4359f728;
  wire al_44b75b16;
  wire al_ab39876a;
  wire al_caca8068;
  wire al_b6bc6cf7;
  wire al_5d326e5d;
  wire al_17c12787;
  wire al_65670e55;
  wire al_15ca3484;
  wire al_e49c184e;
  wire al_c958e833;
  wire al_3e72c22b;
  wire al_12e08f07;
  wire al_65335fa7;
  wire al_df8c0cc2;
  wire al_8e20c85e;
  wire al_2f10c83f;
  wire al_f9924877;
  wire al_26d08bda;
  wire al_e531b722;
  wire al_e8ea4a8d;
  wire al_7d8911c3;
  wire al_4ebe4f9a;
  wire al_a8eab0c8;
  wire al_6567b0f6;
  wire al_72329cb5;
  wire al_c4e45821;
  wire al_aaeb19f7;
  wire al_23e60859;
  wire al_9cb07372;
  wire al_cb712978;
  wire al_7d870001;
  wire al_e748e446;
  wire al_cab235ff;
  wire al_f34da80b;
  wire al_df31c3a1;
  wire al_bb7bf12;
  wire al_1e407f5a;
  wire al_b57079f2;
  wire al_b47584c8;
  wire al_c18c53ba;
  wire al_68105619;
  wire al_386fccc3;
  wire al_cc8bc87f;
  wire al_759d9780;
  wire al_53cc0ecc;
  wire al_2ca2d7bc;
  wire al_f7fcf2a1;
  wire al_fdb8587d;
  wire al_38452a92;
  wire al_b0b78459;
  wire al_6c84cbad;
  wire al_7fa72a5e;
  wire al_59879e6b;
  wire al_41afcc92;
  wire al_b8a226a2;
  wire al_1f6dda96;
  wire al_ae23d17f;
  wire al_86543e7b;
  wire al_2c034ec4;
  wire al_69054c50;
  wire al_3ca382aa;
  wire al_e5156e61;
  wire al_73a263d4;
  wire al_a502ee6;
  wire al_6e5fe692;
  wire al_9fadbc99;
  wire al_7e4e201e;
  wire al_b5f76101;
  wire al_a71f7b3c;
  wire al_6b47e31e;
  wire al_d6e96525;
  wire al_224cbb04;
  wire al_5c961523;
  wire al_146bb661;
  wire al_ae305841;
  wire al_a56ffae1;
  wire al_f5b95ad4;
  wire al_19de37d3;
  wire al_7b57cbb6;
  wire al_4d3e12f0;
  wire al_417e5201;
  wire al_12ccb57b;
  wire al_4e3c3c1e;
  wire al_a68c8fdd;
  wire al_c6b7617c;
  wire al_7ee2af8f;
  wire al_10d4c4b6;
  wire al_aefa880a;
  wire al_dbb207a;
  wire al_94e27914;
  wire al_8abb9d02;
  wire al_420e50cb;
  wire al_42f3bac7;
  wire al_e1983c08;
  wire al_a657a302;
  wire al_46228dd4;
  wire al_d9253b60;
  wire al_9aed2757;
  wire al_ed505fc9;
  wire al_d3c1dd73;
  wire al_b76e4bca;
  wire al_99c75e01;
  wire al_38d9fe9;
  wire al_bd9a895c;
  wire al_13d66540 /* synthesis keep=true */ ;
  wire al_3cc6b708;
  wire al_70117344;
  wire al_9a7b3b80;
  wire al_8cf002a4;
  wire al_b3cfcb5e;
  wire al_f1015bac;
  wire al_fd6a3ba4;
  wire al_42d963e6;
  wire al_4e8fb619;
  wire al_5b144427;
  wire al_142dd1c8;
  wire al_23ce284b;
  wire al_fbdc3092;
  wire al_9929d21;
  wire al_c732c324;
  wire al_ce1c71c5;
  wire al_77d022d8;
  wire al_8815304a;
  wire al_93161d1e;
  wire al_fd460907;
  wire al_e470f61d;
  wire al_5be1fa83;
  wire al_8d08d03c;
  wire al_e2d4d651;
  wire al_8e003744;
  wire al_770f9dd1;
  wire al_d0276689;
  wire al_6e370c03;
  wire al_830e948;
  wire al_25e4ab96;
  wire al_ade031de;
  wire al_7bafa36d;
  wire al_91458dff;
  wire al_8b05cae6;
  wire al_c41fccfb;
  wire al_8dc56974;
  wire al_d2a2bf32;
  wire al_1919cac5;
  wire al_f9c30b23;
  wire al_521fd670;
  wire al_d88aee38;
  wire al_a48594d3;
  wire al_20f5f77c;
  wire al_d27a1279;
  wire al_a771a309;
  wire al_2fc8b96e;
  wire al_eadb4e14;
  wire al_8d8df5a3;
  wire al_1f414bbe;
  wire al_7bbb36d3;
  wire al_4e018b61;
  wire al_6db10ea9;
  wire al_722c0dcd;
  wire al_e2f3bed2;
  wire al_a88d3bd8;
  wire al_24944e5c;
  wire al_3a2d553d;
  wire al_d4c409ba;
  wire al_f9e69b00;
  wire al_4f9aa153;
  wire al_dc57999f;
  wire al_c9d182cf;
  wire al_1f596d24;
  wire al_72ab91cb;
  wire al_7c6973e;
  wire al_df90085e;
  wire al_4ab9f9ad;
  wire al_17b42586;
  wire al_6f07b96e;
  wire al_535f72cd;
  wire al_30c9bd77;
  wire al_843f6bac;
  wire al_1759a3a0;
  wire al_87f40037;
  wire al_e6d4af1;
  wire al_815c8034;
  wire al_8e660235;
  wire al_d90f1fe1;
  wire al_31cf7bc9;
  wire al_10f5be33;
  wire al_be14e3f3;
  wire al_ea6ecc89;
  wire al_335c3c71;
  wire al_8fa72152;
  wire al_fbbf0c04;
  wire al_20c1f74d;
  wire al_b40c9ab5;
  wire al_4aba11ac;
  wire al_ba71435f;
  wire al_2e8aa91;
  wire al_b09b809;
  wire al_6e50ac65;
  wire al_b0c5cb0b;
  wire al_e2476620;
  wire al_ee7571b0;
  wire al_9a6187ef;
  wire al_61d4d1dd;
  wire al_2a05599e;
  wire al_a04a63e0;
  wire al_1a61307;
  wire al_ec12476e;
  wire al_c446e1c1;
  wire al_8ad430a7;
  wire al_9f893f0c;
  wire al_95dd6731;
  wire al_b3610ba2;
  wire al_41f57e5d;
  wire al_dc8a13dc;
  wire al_a0a92d29;
  wire al_70ff6ecf;
  wire al_1c0f25b0;
  wire al_ef98f3e9;
  wire al_d55891ef;
  wire al_92cbdd49;
  wire al_5b5189ed;
  wire al_4f8f3ec;
  wire al_6652ce21;
  wire al_3e851499;
  wire al_c03f902b;
  wire al_787c471e;
  wire al_db74407e;
  wire al_69a4bab5;
  wire al_556566a0;
  wire al_77720e8a;
  wire al_f8edc4ff;
  wire al_925b7c77;
  wire al_4d350d21;
  wire al_db0962eb;
  wire al_cae86888;
  wire al_e5334d53;
  wire al_e0c544fc;
  wire al_6bd0f993;
  wire al_a1041e9;
  wire al_3c6c8ee5;
  wire al_bcb98901;
  wire al_199f1a83;
  wire al_deb7c4e9;
  wire al_1e064d5f;
  wire al_4cc6df6e;
  wire al_ef6225f5;
  wire al_6bddd01a;
  wire al_5f1c8d24;
  wire al_83ebd977;
  wire al_c678f752;
  wire al_c3e70575;
  wire al_3ea78ea2;
  wire al_4864d933;
  wire al_38793d0;
  wire al_4708b339;
  wire al_3ec6ca0b;
  wire al_2efa36ca;
  wire al_e956701b;
  wire al_5e6f3859;
  wire al_d79d15f2;
  wire al_35f768f4;
  wire al_4e23dc54;
  wire al_ee615f87;
  wire al_59fdd957;
  wire al_cc2e5bcc;
  wire al_1bbf8570;
  wire al_31be1d74;
  wire al_14f4e684;
  wire al_b56307ec;
  wire al_2f52bc7e;
  wire al_7cd149c6;
  wire al_652cea26;
  wire al_28d8d34d;
  wire al_89f795c9;
  wire al_a9490be8;
  wire al_8c43abb;
  wire al_9dcab982;
  wire al_46888ef2;
  wire al_2bb74c3d;
  wire al_53b6ba74;
  wire al_80360204;
  wire al_7da0d957;
  wire al_6dc98a03;
  wire al_fa62f20b;
  wire al_df7aa915;
  wire al_49840bbd;
  wire al_796e34c4;
  wire al_74f1ae6b;
  wire al_fef4ecdb;
  wire al_314e2528;
  wire al_b8da0e9e;
  wire al_7ceaf80e;
  wire al_c81182c;
  wire al_fdd1bba3;
  wire al_ab1b2b16;
  wire al_cea991a;
  wire al_64f79045;
  wire al_2c63960b;
  wire al_d9d76d0a;
  wire al_646f260c;
  wire al_3da9562a;
  wire al_8695553e;
  wire al_21d51e65;
  wire al_eda53b41;
  wire al_9f6750b6;
  wire al_860bc871;
  wire al_82133c54;
  wire al_39705b9f;
  wire al_106fddab;
  wire al_33cf56b3;
  wire al_b8cc00cf;
  wire al_228163ab;
  wire al_12b38499;
  wire al_4b7e1c0f;
  wire al_3d66f550;
  wire al_53c183a7;
  wire al_ad58fbc9;
  wire al_b6615be3;
  wire al_ac593c94;
  wire al_c802abc3;
  wire al_f7c9608b;
  wire al_435ecf83;
  wire al_c85cbcb;
  wire al_c600a777;
  wire al_71cac35e;
  wire al_267f05f8;
  wire al_e6ea44e6;
  wire al_55882f9d;
  wire al_9b5a4dbd;
  wire al_26a2c365;
  wire al_4b4a698a;
  wire al_d3da8bb7 /* synthesis keep=true */ ;
  wire al_f5d41495;
  wire al_1342f12a;
  wire al_b00f7d00;
  wire al_411ed67e;
  wire al_7b91dfdd;
  wire al_f4c0ad0d;
  wire al_5d73fdac;
  wire al_d86483c1;
  wire al_4ba727b9;
  wire al_ff9e30e3;
  wire al_62c7fa0b;
  wire al_c77e9fbd;
  wire al_e46ca45e;
  wire al_70f2e5bd;
  wire al_7fe14516;
  wire al_cf62a4e7;
  wire al_2fadb06;
  wire al_cc952326;
  wire al_3cc49650;
  wire al_f567595c;
  wire al_20e796af;
  wire al_710215be;
  wire al_d0805f59;
  wire al_a2b915e0;
  wire al_6c6e8c75;
  wire al_5f044880;
  wire al_1ea20fda;
  wire al_4dade993;
  wire al_d7411c1e;
  wire al_7e6b3b5a;
  wire al_9683b2fb;
  wire al_881adcbc;
  wire al_cb65ad25;
  wire al_b3b929ae;
  wire al_60238e88;
  wire al_2d3877ba;
  wire al_efb91504;
  wire al_2404250b;
  wire al_691fa5a3;
  wire al_37606c32;
  wire al_817a8c80;
  wire al_efea142b;
  wire al_5c1ef4c7;
  wire al_1cb90ce6;
  wire al_ac2df9bf;
  wire al_33994c72;
  wire al_607ca590;
  wire al_e0914439;
  wire al_a28bab3a;
  wire al_4c8ccef5;
  wire al_a390ad74;
  wire al_48ead91e;
  wire al_7d364519;
  wire al_ebd79caa;
  wire al_8f0f91a1;
  wire al_2117afe8;
  wire al_20745547;
  wire al_83931c3d;
  wire al_aa906eb4;
  wire al_72bfbb1a;
  wire al_5f0a94fd;
  wire al_eaa97ed5;
  wire al_54a8a910;
  wire al_f49dc4e0;
  wire al_361b3557;
  wire al_60b9b0f8;
  wire al_41c5883;
  wire al_2acf9590;
  wire al_9c1746a1;
  wire al_f4446f72;
  wire al_9c945a81;
  wire al_a2eb56c3;
  wire al_fb87711d;
  wire al_8c8985a1;
  wire al_99dca23;
  wire al_adc73f46;
  wire al_2db7ae9f;
  wire al_4c1ffe8c;
  wire al_5de748fa;
  wire al_5679c3a4;
  wire al_ba7f7c4;
  wire al_79846c19;
  wire al_42d1f999;
  wire al_c254d68a;
  wire al_2b594476;
  wire al_1dbc8101;
  wire al_1506e6b3;
  wire al_65787e3f;
  wire al_4b87de86;
  wire al_1081a2ca;
  wire al_3d1dbb20;
  wire al_b2e217b;
  wire al_d7967164;
  wire al_c66db911;
  wire al_73668eea;
  wire al_b7e19172;
  wire al_7ab8db7c;
  wire al_994a49f;
  wire al_65ea04b6;
  wire al_4743910a;
  wire al_4fcbf6ef;
  wire al_ddc5d17a;
  wire al_2bfd730a;
  wire al_39c9e6e2;
  wire al_e2323e1d;
  wire al_ce09b21b;
  wire al_73e64072;
  wire al_bd522ea7;
  wire al_792502fb;
  wire al_eefb494d;
  wire al_c0cdd2f2;
  wire al_61b9dbed;
  wire al_e4e2df3a;
  wire al_bd9db94a;
  wire al_2fdd1128;
  wire al_3f1b9f0e;
  wire al_e059f386;
  wire al_54647363;
  wire al_b627b129;
  wire al_31a7d949;
  wire al_fd874a49;
  wire al_7905d584;
  wire al_ba6805c2;
  wire al_957b61e0;
  wire al_9e2fe654;
  wire al_2cac5213;
  wire al_c5c99a19;
  wire al_9b71a4e4;
  wire al_312b2dca;
  wire al_b49bcb3;
  wire al_d8d52ddc;
  wire al_3ed1abca;
  wire al_f07cc0e;
  wire al_a4c76fab;
  wire al_ad24301;
  wire al_8091f068;
  wire al_af74714f;
  wire al_3310bf9b;
  wire al_a6167193;
  wire al_3728ce00;
  wire al_fd1400b6;
  wire al_72450658;
  wire al_733e11d7;
  wire al_2c66a236;
  wire al_e3e65c55;
  wire al_2eb834f5;
  wire al_ec10e78f;
  wire al_e75d67c1;
  wire al_316d230a;
  wire al_6d6f3341;
  wire al_898acbc2;
  wire al_e1d70a3d;
  wire al_fdf8d449;
  wire al_6aad2723;
  wire al_be012e15;
  wire al_3bfb38e8;
  wire al_d2cdc7c9;
  wire al_84ac14c0;
  wire al_1b504c84;
  wire al_a6be8738;
  wire al_c21b49ee;
  wire al_b09bcab2;
  wire al_b62a0a78;
  wire al_27d43db3;
  wire al_d9a683f3;
  wire al_7aee3607;
  wire al_852588b2;
  wire al_664e4e8f;
  wire al_6f9c4eba;
  wire al_55b9d73d;
  wire al_3858b210;
  wire al_96b7453;
  wire al_ee3904b1;
  wire al_1abf75fc;
  wire al_f9fd3044;
  wire al_14656fdb;
  wire al_cda79e31;
  wire al_130738c8;
  wire al_f45ad02a;
  wire al_4783da3f;
  wire al_b285e414;
  wire al_ef6d9f73;
  wire al_a7a585be;
  wire al_3f68feff;
  wire al_92250858;
  wire al_b4d25a49;
  wire al_3b280eeb;
  wire al_e3bba389;
  wire al_a07095e8;
  wire al_bf50c51c;
  wire al_472a7b46;
  wire al_b9b495b9;
  wire al_4531bc64;
  wire al_3f7b50be;
  wire al_4cb605a3;
  wire al_2ebef479;
  wire al_d93c50d7;
  wire al_6a0200a0;
  wire al_15554a76;
  wire al_ce868614;
  wire al_89b57934;
  wire al_d6502391;
  wire al_b57594f0;
  wire al_ca5b293f;
  wire al_da329b96;
  wire al_f3b50940;
  wire al_14200974;
  wire al_71fc1ad7;
  wire al_6db5b9d2;
  wire al_b8212fd4;
  wire al_1584b2ff;
  wire al_e463a453;
  wire al_952b0ccf;
  wire al_bf72b0fb;
  wire al_221290fc;
  wire al_fd118264;
  wire al_f3b3330;
  wire al_6adcd3f0;
  wire al_dd36eaa4;
  wire al_7c446883;
  wire al_86df7d12;
  wire al_1591047a;
  wire al_d3c4d360;
  wire al_6d6760dd;
  wire al_9cf6a965;
  wire al_37a8c4a3;
  wire al_2c31bcd7;
  wire al_bbe31482;
  wire al_edff11e6;
  wire al_4b287773;
  wire al_a18a78ec;
  wire al_f8b11b95;
  wire al_dd0c66b3;
  wire al_edb83574;
  wire al_2935d0ed;
  wire al_538eda90;
  wire al_2503fdb;
  wire al_f8fcd204;
  wire al_467a2ca;
  wire al_c76ae5c3;
  wire al_d2c8f1b1;
  wire al_282d371d;
  wire al_cd27f05c;
  wire al_27b77d58;
  wire al_d4d145cc;
  wire al_129a2529;
  wire al_14cefac2;
  wire al_6fd6ffff;
  wire al_f645b571;
  wire al_3419432c;
  wire al_b9e4ee74;
  wire al_4b747cba;
  wire al_733c48ff;
  wire al_5e87f1a6;
  wire al_addcc22;
  wire al_549369e;
  wire al_e837a56c;
  wire al_3021b8d9;
  wire al_984d7f7;
  wire al_f24aaa07;
  wire al_f9e997a5;
  wire al_1819221f;
  wire al_555b330b;
  wire al_44a10d10;
  wire al_555cabbf;
  wire al_8f3c4595;
  wire al_3daf893a /* synthesis keep=true */ ;
  wire al_6ab6f142;
  wire al_947c0ab9;
  wire al_2b896d2b /* synthesis keep=true */ ;
  wire al_e6043332;
  wire al_6d2ef296 /* synthesis keep=true */ ;
  wire al_9431cde9;
  wire al_4fdebbe9 /* synthesis keep=true */ ;
  wire al_b456bf15;
  wire al_d56bc9f8 /* synthesis keep=true */ ;
  wire al_fd258f8;
  wire al_630d6511 /* synthesis keep=true */ ;
  wire al_1ceb77fa;
  wire al_ba561a9e /* synthesis keep=true */ ;
  wire al_d872bb7e;
  wire al_64b5f594 /* synthesis keep=true */ ;
  wire al_b9b87e33;
  wire al_3730b5bd;
  wire al_e4f5976f /* synthesis keep=true */ ;
  wire al_2ca0cac1;
  wire al_a36f4fe4;
  wire al_e0470675;
  wire al_1c2bc502;
  wire al_fba0e4a3;
  wire al_8a002c3c;
  wire al_9056b393;
  wire al_44ed9c4;
  wire al_a33220fb;
  wire al_78b4c22e;
  wire al_55e87168;
  wire al_1fc0eb8a;
  wire al_5e51060a;
  wire al_aa3cad87;
  wire al_33ae520;
  wire al_9a26ce4f;
  wire al_b8363901;
  wire al_603c814;
  wire al_6b7d1c4;
  wire al_5ed629c8;
  wire al_2d1611fb;
  wire al_6c6fd169;
  wire al_7bc48670;
  wire al_b03fffe1;
  wire al_cf2346e1;
  wire al_d22a1e42;
  wire al_17f22329;

  assign al_ef3696df[0] = clk;
  assign ddr_app_wdf_rdy = al_6ab6f142;
  assign dfi_act_n_p[3] = dfi_act_n_p[0];
  assign dfi_act_n_p[2] = dfi_act_n_p[0];
  assign dfi_address_p[55] = dfi_address_p[42];
  assign dfi_address_p[54] = dfi_address_p[42];
  assign dfi_address_p[53] = dfi_address_p[42];
  assign dfi_address_p[52] = dfi_address_p[42];
  assign dfi_address_p[51] = dfi_address_p[42];
  assign dfi_address_p[50] = dfi_address_p[42];
  assign dfi_address_p[49] = dfi_address_p[42];
  assign dfi_address_p[48] = dfi_address_p[42];
  assign dfi_address_p[47] = dfi_address_p[42];
  assign dfi_address_p[46] = dfi_address_p[42];
  assign dfi_address_p[45] = dfi_address_p[42];
  assign dfi_address_p[44] = dfi_address_p[42];
  assign dfi_address_p[43] = dfi_address_p[42];
  assign dfi_address_p[41] = 1'b0;
  assign dfi_address_p[40] = 1'b0;
  assign dfi_address_p[39] = 1'b0;
  assign dfi_address_p[38] = 1'b0;
  assign dfi_address_p[37] = 1'b0;
  assign dfi_address_p[36] = 1'b0;
  assign dfi_address_p[35] = 1'b0;
  assign dfi_address_p[34] = 1'b0;
  assign dfi_address_p[33] = 1'b0;
  assign dfi_address_p[32] = 1'b0;
  assign dfi_address_p[31] = 1'b0;
  assign dfi_address_p[30] = 1'b0;
  assign dfi_address_p[29] = 1'b0;
  assign dfi_address_p[28] = 1'b0;
  assign dfi_address_p[13] = 1'b0;
  assign dfi_address_p[12] = 1'b0;
  assign dfi_address_p[11] = 1'b0;
  assign dfi_address_p[10] = 1'b0;
  assign dfi_address_p[2] = 1'b0;
  assign dfi_address_p[1] = 1'b0;
  assign dfi_bank_p[8] = 1'b0;
  assign dfi_bank_p[7] = 1'b0;
  assign dfi_bank_p[6] = 1'b0;
  assign dfi_cas_n_p[2] = dfi_act_n_p[0];
  assign dfi_cas_n_p[1] = dfi_act_n_p[0];
  assign dfi_cke_p[2] = dfi_cke_p[0];
  assign dfi_cke_p[1] = dfi_cke_p[0];
  assign dfi_cs_n_p[2] = dfi_act_n_p[0];
  assign dfi_cs_n_p[1] = dfi_act_n_p[1];
  assign dfi_cs_n_p[0] = dfi_cas_n_p[0];
  assign dfi_odt_p[3] = dfi_odt_p[2];
  assign dfi_odt_p[1] = dfi_odt_p[0];
  assign dfi_ras_n_p[2] = dfi_act_n_p[0];
  assign dfi_ras_n_p[1] = dfi_act_n_p[1];
  assign dfi_ras_n_p[0] = dfi_act_n_p[0];
  assign dfi_rddata_en_p[15] = dfi_rddata_en_p[12];
  assign dfi_rddata_en_p[14] = dfi_rddata_en_p[12];
  assign dfi_rddata_en_p[13] = dfi_rddata_en_p[12];
  assign dfi_rddata_en_p[11] = dfi_rddata_en_p[8];
  assign dfi_rddata_en_p[10] = dfi_rddata_en_p[8];
  assign dfi_rddata_en_p[9] = dfi_rddata_en_p[8];
  assign dfi_rddata_en_p[7] = dfi_rddata_en_p[0];
  assign dfi_rddata_en_p[6] = dfi_rddata_en_p[0];
  assign dfi_rddata_en_p[5] = dfi_rddata_en_p[0];
  assign dfi_rddata_en_p[4] = dfi_rddata_en_p[0];
  assign dfi_rddata_en_p[3] = dfi_rddata_en_p[0];
  assign dfi_rddata_en_p[2] = dfi_rddata_en_p[0];
  assign dfi_rddata_en_p[1] = dfi_rddata_en_p[0];
  assign dfi_reset_n[3] = 1'b1;
  assign dfi_reset_n[2] = 1'b1;
  assign dfi_reset_n[1] = 1'b1;
  assign dfi_reset_n[0] = 1'b1;
  assign dfi_we_n_p[2] = dfi_act_n_p[0];
  assign dfi_we_n_p[1] = dfi_act_n_p[0];
  assign dfi_wrdata_en_p[15] = dfi_wrdata_en_p[12];
  assign dfi_wrdata_en_p[14] = dfi_wrdata_en_p[12];
  assign dfi_wrdata_en_p[13] = dfi_wrdata_en_p[12];
  assign dfi_wrdata_en_p[11] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[10] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[9] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[8] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[7] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[6] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[5] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[4] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[3] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[2] = dfi_wrdata_en_p[0];
  assign dfi_wrdata_en_p[1] = dfi_wrdata_en_p[0];
  AL_MAP_LUT6 #(
    .EQN("(F*~(~(~E*D*~C)*~(~B*~A)))"),
    .INIT(64'h11111f1100000000))
    al_81464152 (
    .a(al_4732ba15[0]),
    .b(al_4732ba15[1]),
    .c(al_72785055[0]),
    .d(al_72785055[2]),
    .e(al_72785055[1]),
    .f(al_cc4d831c[0]),
    .o(al_80aa352a));
  AL_DFF_0 al_78220107 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9120ce24),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f9840a37));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_1bdfb83a (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_f62f60e1[0]),
    .d(al_7b737f75[0]),
    .e(al_d7fecbad[0]),
    .f(al_8d302088[0]),
    .o(al_9e51440f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_958c2db3 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_cdd95abd[0]),
    .d(al_c5d3b031[0]),
    .e(al_79af3182[0]),
    .f(al_efab6074[0]),
    .o(al_3235c6b2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h333355550f0f00ff))
    al_e6c52c5b (
    .a(al_d81bfd7d),
    .b(al_f3aabbcb),
    .c(al_8d9f1a8e),
    .d(al_3235c6b2),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_f6ab792b));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    al_328d5254 (
    .a(al_4030306c),
    .b(al_f6ab792b),
    .c(al_d1b0929d),
    .d(al_194afe0a[4]),
    .o(al_71c87c87[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_edf785c1 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_41bdf331[0]),
    .d(al_9d72d808[0]),
    .e(al_905e5060[0]),
    .f(al_62b22b32[0]),
    .o(al_12509175));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_565794db (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_af419986[0]),
    .d(al_cf0afe9a[0]),
    .e(al_f594a8d9[0]),
    .f(al_df5cbc72[0]),
    .o(al_3a6224d6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_45886bcc (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_95e9fdd1[0]),
    .d(al_84027ae7[0]),
    .e(al_9f61035a[0]),
    .f(al_4e28198f[0]),
    .o(al_b7e8ef76));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_794f93fb (
    .a(al_9e51440f),
    .b(al_12509175),
    .c(al_3a6224d6),
    .d(al_b7e8ef76),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_4030306c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_23d8e2e (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_74387eee[0]),
    .d(al_c7b20b0[0]),
    .e(al_ff281ad1[0]),
    .f(al_effd30c4[0]),
    .o(al_d81bfd7d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_1141103f (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_adfe279[0]),
    .d(al_eec6554e[0]),
    .e(al_c58c2706[0]),
    .f(al_b1296b3[0]),
    .o(al_f3aabbcb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_f49f9b79 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_a6fdde80[0]),
    .d(al_e6b17901[0]),
    .e(al_57e2199e[0]),
    .f(al_48ac75ce[0]),
    .o(al_8d9f1a8e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_2ccfb3c (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_f62f60e1[1]),
    .d(al_7b737f75[1]),
    .e(al_d7fecbad[1]),
    .f(al_8d302088[1]),
    .o(al_cff749bd));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_18d7ddd7 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_74387eee[1]),
    .d(al_c7b20b0[1]),
    .e(al_ff281ad1[1]),
    .f(al_effd30c4[1]),
    .o(al_cd1bc23c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_693c90db (
    .a(al_e65434a9),
    .b(al_955d2d0b),
    .c(al_761b87c7),
    .d(al_cd1bc23c),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_d3acc8ad));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    al_a60ffe3a (
    .a(al_10c16c),
    .b(al_d3acc8ad),
    .c(al_d1b0929d),
    .d(al_194afe0a[4]),
    .o(al_71c87c87[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_dbb73d40 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_41bdf331[1]),
    .d(al_9d72d808[1]),
    .e(al_905e5060[1]),
    .f(al_62b22b32[1]),
    .o(al_83946844));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_bcaaf242 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_af419986[1]),
    .d(al_cf0afe9a[1]),
    .e(al_f594a8d9[1]),
    .f(al_df5cbc72[1]),
    .o(al_638fd104));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_7308d2cd (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_95e9fdd1[1]),
    .d(al_84027ae7[1]),
    .e(al_9f61035a[1]),
    .f(al_4e28198f[1]),
    .o(al_4edaac38));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_6101f7c7 (
    .a(al_cff749bd),
    .b(al_83946844),
    .c(al_638fd104),
    .d(al_4edaac38),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_10c16c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_6cf913c6 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_a6fdde80[1]),
    .d(al_e6b17901[1]),
    .e(al_57e2199e[1]),
    .f(al_48ac75ce[1]),
    .o(al_e65434a9));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_a4672331 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_cdd95abd[1]),
    .d(al_c5d3b031[1]),
    .e(al_79af3182[1]),
    .f(al_efab6074[1]),
    .o(al_955d2d0b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_7c903dc4 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_adfe279[1]),
    .d(al_eec6554e[1]),
    .e(al_c58c2706[1]),
    .f(al_b1296b3[1]),
    .o(al_761b87c7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_c3fa778a (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_f62f60e1[2]),
    .d(al_7b737f75[2]),
    .e(al_d7fecbad[2]),
    .f(al_8d302088[2]),
    .o(al_8370ebfb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_1cc4dd3b (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_cdd95abd[2]),
    .d(al_c5d3b031[2]),
    .e(al_79af3182[2]),
    .f(al_efab6074[2]),
    .o(al_b7f132ea));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h333355550f0f00ff))
    al_a1245743 (
    .a(al_8c295dd7),
    .b(al_fdbc6cb0),
    .c(al_33827427),
    .d(al_b7f132ea),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_34945d75));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    al_6500682c (
    .a(al_8abdf99c),
    .b(al_34945d75),
    .c(al_d1b0929d),
    .d(al_194afe0a[4]),
    .o(al_71c87c87[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_87fe66bb (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_41bdf331[2]),
    .d(al_9d72d808[2]),
    .e(al_905e5060[2]),
    .f(al_62b22b32[2]),
    .o(al_62f041ec));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_c9bf84f1 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_af419986[2]),
    .d(al_cf0afe9a[2]),
    .e(al_f594a8d9[2]),
    .f(al_df5cbc72[2]),
    .o(al_62b064bd));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_dea77898 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_95e9fdd1[2]),
    .d(al_84027ae7[2]),
    .e(al_9f61035a[2]),
    .f(al_4e28198f[2]),
    .o(al_e5820766));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_cf81a19d (
    .a(al_8370ebfb),
    .b(al_62f041ec),
    .c(al_62b064bd),
    .d(al_e5820766),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_8abdf99c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_d543cf29 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_74387eee[2]),
    .d(al_c7b20b0[2]),
    .e(al_ff281ad1[2]),
    .f(al_effd30c4[2]),
    .o(al_8c295dd7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_bd54695f (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_adfe279[2]),
    .d(al_eec6554e[2]),
    .e(al_c58c2706[2]),
    .f(al_b1296b3[2]),
    .o(al_fdbc6cb0));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_4bbb554a (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_a6fdde80[2]),
    .d(al_e6b17901[2]),
    .e(al_57e2199e[2]),
    .f(al_48ac75ce[2]),
    .o(al_33827427));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_b742390d (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_f62f60e1[3]),
    .d(al_7b737f75[3]),
    .e(al_d7fecbad[3]),
    .f(al_8d302088[3]),
    .o(al_2f53f65));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_22251bbc (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_74387eee[3]),
    .d(al_c7b20b0[3]),
    .e(al_ff281ad1[3]),
    .f(al_effd30c4[3]),
    .o(al_ddf7a9aa));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_7baad471 (
    .a(al_3e22da4d),
    .b(al_b030bf9a),
    .c(al_c2f4eaf6),
    .d(al_ddf7a9aa),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_ef1fe31d));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    al_568b7246 (
    .a(al_b8516693),
    .b(al_ef1fe31d),
    .c(al_d1b0929d),
    .d(al_194afe0a[4]),
    .o(al_71c87c87[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_fce5249a (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_41bdf331[3]),
    .d(al_9d72d808[3]),
    .e(al_905e5060[3]),
    .f(al_62b22b32[3]),
    .o(al_d0d67001));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_773bdfc (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_af419986[3]),
    .d(al_cf0afe9a[3]),
    .e(al_f594a8d9[3]),
    .f(al_df5cbc72[3]),
    .o(al_a7c3fab2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_c1ca3934 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_95e9fdd1[3]),
    .d(al_84027ae7[3]),
    .e(al_9f61035a[3]),
    .f(al_4e28198f[3]),
    .o(al_505af09f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_273f0e15 (
    .a(al_2f53f65),
    .b(al_d0d67001),
    .c(al_a7c3fab2),
    .d(al_505af09f),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_b8516693));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_d11a39cc (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_a6fdde80[3]),
    .d(al_e6b17901[3]),
    .e(al_57e2199e[3]),
    .f(al_48ac75ce[3]),
    .o(al_3e22da4d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_5e9d1eb8 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_cdd95abd[3]),
    .d(al_c5d3b031[3]),
    .e(al_79af3182[3]),
    .f(al_efab6074[3]),
    .o(al_b030bf9a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_efafa617 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_adfe279[3]),
    .d(al_eec6554e[3]),
    .e(al_c58c2706[3]),
    .f(al_b1296b3[3]),
    .o(al_c2f4eaf6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_db5298ea (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_95e9fdd1[4]),
    .d(al_84027ae7[4]),
    .e(al_9f61035a[4]),
    .f(al_4e28198f[4]),
    .o(al_6bbf1231));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_716918ae (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_74387eee[4]),
    .d(al_c7b20b0[4]),
    .e(al_ff281ad1[4]),
    .f(al_effd30c4[4]),
    .o(al_35f5fbe2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_e3675b33 (
    .a(al_5cfcbe8d),
    .b(al_78f859ca),
    .c(al_9cac2c36),
    .d(al_35f5fbe2),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_37d972e0));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    al_188b4a34 (
    .a(al_a87038a),
    .b(al_37d972e0),
    .c(al_d1b0929d),
    .d(al_194afe0a[4]),
    .o(al_71c87c87[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_de0ed7ba (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_af419986[4]),
    .d(al_cf0afe9a[4]),
    .e(al_f594a8d9[4]),
    .f(al_df5cbc72[4]),
    .o(al_2b0ac92a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_f2fe0443 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_f62f60e1[4]),
    .d(al_7b737f75[4]),
    .e(al_d7fecbad[4]),
    .f(al_8d302088[4]),
    .o(al_f9950e01));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_6f3ac160 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_41bdf331[4]),
    .d(al_9d72d808[4]),
    .e(al_905e5060[4]),
    .f(al_62b22b32[4]),
    .o(al_f4c5dfba));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h333355550f0f00ff))
    al_6a4155af (
    .a(al_6bbf1231),
    .b(al_2b0ac92a),
    .c(al_f9950e01),
    .d(al_f4c5dfba),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_a87038a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_cbbda4e4 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_a6fdde80[4]),
    .d(al_e6b17901[4]),
    .e(al_57e2199e[4]),
    .f(al_48ac75ce[4]),
    .o(al_5cfcbe8d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_ba04107e (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_cdd95abd[4]),
    .d(al_c5d3b031[4]),
    .e(al_79af3182[4]),
    .f(al_efab6074[4]),
    .o(al_78f859ca));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_dd19d2f (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_adfe279[4]),
    .d(al_eec6554e[4]),
    .e(al_c58c2706[4]),
    .f(al_b1296b3[4]),
    .o(al_9cac2c36));
  AL_DFF_0 al_ac407fa7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d1b0929d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9841dcd3));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_45865a0c (
    .a(dfi_rddata_valid_w[15]),
    .b(dfi_rddata_valid_w[14]),
    .c(dfi_rddata_valid_w[13]),
    .d(dfi_rddata_valid_w[12]),
    .o(al_c6c76177));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_c49929e9 (
    .a(dfi_rddata_valid_w[7]),
    .b(dfi_rddata_valid_w[6]),
    .c(dfi_rddata_valid_w[5]),
    .d(dfi_rddata_valid_w[4]),
    .o(al_95b46020));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_5cbd16a0 (
    .a(al_95b46020),
    .b(dfi_rddata_valid_w[3]),
    .c(dfi_rddata_valid_w[2]),
    .d(dfi_rddata_valid_w[1]),
    .e(dfi_rddata_valid_w[0]),
    .o(al_95467c49));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~E*~D*~C*B*A)"),
    .INIT(64'hfffffffffffffff7))
    al_908ffe3e (
    .a(al_95467c49),
    .b(al_c6c76177),
    .c(dfi_rddata_valid_w[11]),
    .d(dfi_rddata_valid_w[10]),
    .e(dfi_rddata_valid_w[9]),
    .f(dfi_rddata_valid_w[8]),
    .o(al_4779567c));
  AL_DFF_0 al_f1170662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4779567c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1b0929d));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(~C*B*A))"),
    .INIT(16'hff08))
    al_5b1b1a35 (
    .a(al_f9840a37),
    .b(al_4732ba15[0]),
    .c(al_4732ba15[1]),
    .d(al_c0f3a3cd[7]),
    .o(al_4aabc590[0]));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*A*~(~C*B))"),
    .INIT(64'h00000000a2000000))
    al_7ee1e69a (
    .a(al_f9840a37),
    .b(al_4732ba15[0]),
    .c(al_4732ba15[1]),
    .d(al_72785055[0]),
    .e(al_72785055[2]),
    .f(al_72785055[1]),
    .o(al_4aabc590[4]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(~D*C*B))"),
    .INIT(16'haaea))
    al_fedd6419 (
    .a(al_4aabc590[4]),
    .b(al_f9840a37),
    .c(al_4732ba15[0]),
    .d(al_4732ba15[1]),
    .o(al_4aabc590[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_594e1ff9 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_f62f60e1[5]),
    .d(al_7b737f75[5]),
    .e(al_d7fecbad[5]),
    .f(al_8d302088[5]),
    .o(al_d31b0b8f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_d9b9026b (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_74387eee[5]),
    .d(al_c7b20b0[5]),
    .e(al_ff281ad1[5]),
    .f(al_effd30c4[5]),
    .o(al_6051bc62));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_2f8809f2 (
    .a(al_96b41fb2),
    .b(al_cc069a1e),
    .c(al_66f9507b),
    .d(al_6051bc62),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_48c4d402));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    al_320a1146 (
    .a(al_24ea9f76),
    .b(al_48c4d402),
    .c(al_d1b0929d),
    .d(al_194afe0a[4]),
    .o(al_e3d7dc13));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_7533dc7b (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_41bdf331[5]),
    .d(al_9d72d808[5]),
    .e(al_905e5060[5]),
    .f(al_62b22b32[5]),
    .o(al_8f66e49d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_5b9b7336 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_af419986[5]),
    .d(al_cf0afe9a[5]),
    .e(al_f594a8d9[5]),
    .f(al_df5cbc72[5]),
    .o(al_20ccc531));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_a49a27d0 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_95e9fdd1[5]),
    .d(al_84027ae7[5]),
    .e(al_9f61035a[5]),
    .f(al_4e28198f[5]),
    .o(al_eac4076b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff55553333))
    al_4939bbcd (
    .a(al_d31b0b8f),
    .b(al_8f66e49d),
    .c(al_20ccc531),
    .d(al_eac4076b),
    .e(al_194afe0a[2]),
    .f(al_194afe0a[3]),
    .o(al_24ea9f76));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_45c81099 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_a6fdde80[5]),
    .d(al_e6b17901[5]),
    .e(al_57e2199e[5]),
    .f(al_48ac75ce[5]),
    .o(al_96b41fb2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_4099f76c (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_cdd95abd[5]),
    .d(al_c5d3b031[5]),
    .e(al_79af3182[5]),
    .f(al_efab6074[5]),
    .o(al_cc069a1e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_75df8869 (
    .a(al_194afe0a[0]),
    .b(al_194afe0a[1]),
    .c(al_adfe279[5]),
    .d(al_eec6554e[5]),
    .e(al_c58c2706[5]),
    .f(al_b1296b3[5]),
    .o(al_66f9507b));
  AL_DFF_0 al_42ce5c6f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3d7dc13),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7a04bdba));
  AL_DFF_0 al_202ace5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44c9e0a6[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_act_n_p[0]));
  AL_DFF_0 al_213526da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e84b9bda[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_act_n_p[1]));
  AL_DFF_0 al_9cf9c1ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44c9e0a6[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_cas_n_p[0]));
  AL_DFF_0 al_d4158be3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44c9e0a6[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_cas_n_p[3]));
  AL_DFF_0 al_494f86ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33061d84[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44c9e0a6[0]));
  AL_DFF_0 al_8f13272f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33061d84[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44c9e0a6[1]));
  AL_DFF_0 al_eeba1c6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33061d84[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44c9e0a6[3]));
  AL_DFF_0 al_7e35553a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a4f25695),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33061d84[0]));
  AL_DFF_0 al_cec6b81 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(1'b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33061d84[1]));
  AL_DFF_0 al_221e893c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97dc1b67),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33061d84[3]));
  AL_DFF_0 al_796d084b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2cf67988[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_cke_p[0]));
  AL_DFF_0 al_594f7ed7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2cf67988[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_cke_p[3]));
  AL_DFF_0 al_77958966 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55586ac1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2cf67988[0]));
  AL_DFF_0 al_9c7333e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55586ac1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2cf67988[3]));
  AL_DFF_0 al_5cc55830 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_45d6e796[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55586ac1[0]));
  AL_DFF_0 al_adb79c2e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff1cf72f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55586ac1[3]));
  AL_DFF_0 al_566511d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e84b9bda[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_cs_n_p[3]));
  AL_DFF_0 al_a86de90a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ac432c54[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e84b9bda[1]));
  AL_DFF_0 al_a6a5d6ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ac432c54[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e84b9bda[3]));
  AL_DFF_0 al_e63f26ff (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56820b3e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac432c54[1]));
  AL_DFF_0 al_16fcc833 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56820b3e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac432c54[3]));
  AL_DFF_0 al_2062ebb6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_49010dd2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_odt_p[0]));
  AL_DFF_0 al_d1141260 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_49010dd2[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_odt_p[2]));
  AL_DFF_0 al_cd5ee54d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5dbfdac[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49010dd2[0]));
  AL_DFF_0 al_91b2301d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5dbfdac[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49010dd2[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d70afa99 (
    .a(al_be11f694),
    .b(al_ef9accde),
    .o(al_16ace516[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_4742273a (
    .a(al_16ace516[27]),
    .b(rst),
    .c(al_e5dbfdac[2]),
    .o(al_159f33b5));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .INIT(16'hf3e2))
    al_f70f05de (
    .a(al_16ace516[27]),
    .b(rst),
    .c(al_e5dbfdac[0]),
    .d(al_dc65c0d1[21]),
    .o(al_86a56c9a));
  AL_DFF_0 al_70e0f5ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_86a56c9a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e5dbfdac[0]));
  AL_DFF_0 al_2c7822b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_159f33b5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e5dbfdac[2]));
  AL_DFF_0 al_510ebef8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_733ec639[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_ras_n_p[3]));
  AL_DFF_0 al_ddae5c1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3d66861c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_733ec639[3]));
  AL_DFF_0 al_a3517000 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6c456f4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d66861c[3]));
  AL_DFF_0 al_5183ec50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0f3a3cd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_rddata_en_p[0]));
  AL_DFF_0 al_736a8853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0f3a3cd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_rddata_en_p[8]));
  AL_DFF_0 al_db8e87fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0f3a3cd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_rddata_en_p[12]));
  AL_DFF_0 al_508c239a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_94b2715c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_we_n_p[0]));
  AL_DFF_0 al_b07bf5a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_94b2715c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_we_n_p[3]));
  AL_DFF_0 al_412f0729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b99d9508[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_94b2715c[0]));
  AL_DFF_0 al_20646ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b99d9508[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_94b2715c[3]));
  AL_DFF_0 al_3061cdb7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1dd73244),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b99d9508[0]));
  AL_DFF_0 al_13061730 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2ccfdf18),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b99d9508[3]));
  AL_DFF_0 al_dbb221a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8679dfa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_en_p[0]));
  AL_DFF_0 al_be3cf266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8679dfa[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_en_p[12]));
  AL_DFF_0 al_5993376c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4732ba15[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4732ba15[3]));
  AL_DFF_0 al_43a3f556 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4732ba15[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4732ba15[4]));
  AL_DFF_0 al_3a7269e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4732ba15[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4da789e[0]));
  AL_DFF_0 al_e1186f9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4732ba15[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4da789e[1]));
  AL_DFF_1 al_2816e367 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1dd73244),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4732ba15[0]));
  AL_DFF_1 al_3029ee5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a4f25695),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4732ba15[1]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_bfcb93d5 (
    .a(al_16ace516[27]),
    .o(al_1dd73244));
  AL_DFF_0 al_1e381bc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(1'b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2a9196a6[3]));
  AL_DFF_0 al_32a4d383 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2a9196a6[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48eb6d34[0]));
  AL_DFF_0 al_4419bdf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2ccfdf18),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_72785055[0]));
  AL_DFF_0 al_151b7161 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6c456f4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_72785055[2]));
  AL_DFF_0 al_d2cbb898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_72785055[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_72785055[3]));
  AL_DFF_0 al_dcb4e0ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_72785055[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_72785055[4]));
  AL_DFF_0 al_9102257b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_72785055[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_72785055[5]));
  AL_DFF_0 al_ad176d74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_72785055[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9b4cc10[0]));
  AL_DFF_0 al_824155ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_72785055[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9b4cc10[1]));
  AL_DFF_0 al_c6abe589 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_72785055[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9b4cc10[2]));
  AL_DFF_1 al_42849273 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97dc1b67),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_72785055[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_d09309e4 (
    .a(al_90a0fe97[0]),
    .b(al_8932a489),
    .c(al_165f2734),
    .d(al_4c58e022),
    .o(al_46b8ac3c));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*~(~C*~(E*~D))))"),
    .INIT(32'h2a222a2a))
    al_abdccb5d (
    .a(al_46b8ac3c),
    .b(al_4ba8484b),
    .c(al_4f7a36e8),
    .d(al_c5705f8a),
    .e(al_11b28491),
    .o(al_2ccfdf18));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    al_3522f810 (
    .a(al_46b8ac3c),
    .b(al_4ba8484b),
    .c(al_4f7a36e8),
    .d(al_c5705f8a),
    .o(al_e6c456f4));
  AL_MAP_LUT4 #(
    .EQN("~(D*~C*B*A)"),
    .INIT(16'hf7ff))
    al_5c9a779b (
    .a(al_46b8ac3c),
    .b(al_4ba8484b),
    .c(al_4f7a36e8),
    .d(al_c5705f8a),
    .o(al_97dc1b67));
  AL_DFF_0 al_6300fe06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[0]));
  AL_DFF_0 al_f6dbd28a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[3]));
  AL_DFF_0 al_824ee760 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[4]));
  AL_DFF_0 al_9f411b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[5]));
  AL_DFF_0 al_67e3c4c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[6]));
  AL_DFF_0 al_64c39b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[7]));
  AL_DFF_0 al_975e4f61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[8]));
  AL_DFF_0 al_f0ab98e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[9]));
  AL_DFF_0 al_a6a99dd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[14]));
  AL_DFF_0 al_aa7ff3c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[15]));
  AL_DFF_0 al_c8aec549 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[16]));
  AL_DFF_0 al_63698251 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[17]));
  AL_DFF_0 al_66216df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[18]));
  AL_DFF_0 al_a87981a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[19]));
  AL_DFF_0 al_89bb185f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[20]));
  AL_DFF_0 al_7157c4cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[21]));
  AL_DFF_0 al_c81f4fc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[22]));
  AL_DFF_0 al_2e3bfb44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[23]));
  AL_DFF_0 al_896a2fdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[24]));
  AL_DFF_0 al_434d2658 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[25]));
  AL_DFF_0 al_8af830a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[26]));
  AL_DFF_0 al_6280aeb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[27]));
  AL_DFF_0 al_c577d3bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f09d84cf[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_address_p[42]));
  AL_DFF_0 al_c0826e47 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_31c39442),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_194afe0a[3]));
  AL_DFF_0 al_947481d0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c9e6a24c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_194afe0a[4]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_59b82114 (
    .a(al_d1b0929d),
    .b(al_194afe0a[0]),
    .o(al_445ee5b3));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    al_1f952364 (
    .a(al_d1b0929d),
    .b(al_194afe0a[0]),
    .c(al_194afe0a[1]),
    .o(al_44ab4bb8));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*A))"),
    .INIT(16'h7f80))
    al_cf492fac (
    .a(al_d1b0929d),
    .b(al_194afe0a[0]),
    .c(al_194afe0a[1]),
    .d(al_194afe0a[2]),
    .o(al_85b0e5ae));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*C*B*A))"),
    .INIT(32'h7fff8000))
    al_40dc885e (
    .a(al_d1b0929d),
    .b(al_194afe0a[0]),
    .c(al_194afe0a[1]),
    .d(al_194afe0a[2]),
    .e(al_194afe0a[3]),
    .o(al_31c39442));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_687440ef (
    .a(al_d1b0929d),
    .b(al_194afe0a[0]),
    .c(al_194afe0a[1]),
    .d(al_194afe0a[2]),
    .e(al_194afe0a[3]),
    .f(al_194afe0a[4]),
    .o(al_c9e6a24c));
  AL_DFF_0 al_cb42d9a7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_445ee5b3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_194afe0a[0]));
  AL_DFF_0 al_a8b6fa46 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44ab4bb8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_194afe0a[1]));
  AL_DFF_0 al_8140a772 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_85b0e5ae),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_194afe0a[2]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_6f73e438 (
    .a(al_643bfe7d),
    .b(al_950c19d6),
    .c(al_efab6074[3]),
    .o(al_776135fb));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_879d469 (
    .a(al_950c19d6),
    .b(al_efab6074[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_4c1ceb3d));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*C*~B*A)"),
    .INIT(64'h0000200000000000))
    al_28872c82 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_e0ba4c33));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a6638a18 (
    .a(al_95c3862c),
    .b(al_e0ba4c33),
    .c(al_57e2199e[4]),
    .o(al_7ebd1ee0));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_6e3009ce (
    .a(al_5083706f),
    .b(al_e0ba4c33),
    .c(al_57e2199e[0]),
    .o(al_462dcba0));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_b6488c13 (
    .a(al_f6411514),
    .b(al_e0ba4c33),
    .c(al_57e2199e[1]),
    .o(al_13f4f154));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_675fa34c (
    .a(al_6f628420),
    .b(al_e0ba4c33),
    .c(al_57e2199e[2]),
    .o(al_1ec9bae4));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_4d1e2063 (
    .a(al_643bfe7d),
    .b(al_e0ba4c33),
    .c(al_57e2199e[3]),
    .o(al_b87141aa));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_50d6395a (
    .a(al_e0ba4c33),
    .b(al_57e2199e[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_d735f43c));
  AL_DFF_0 al_ebe8abfa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b6e3903),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41bdf331[0]));
  AL_DFF_0 al_4d90dcda (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f32b3ce),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41bdf331[1]));
  AL_DFF_0 al_55ea06c9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a3ec7d2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41bdf331[2]));
  AL_DFF_0 al_ab208fde (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1867b14e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41bdf331[3]));
  AL_DFF_0 al_faa3a1b1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_595cd185),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41bdf331[4]));
  AL_DFF_0 al_77fa7ff4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d5c31119),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41bdf331[5]));
  AL_DFF_0 al_60425702 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dc426867),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d72d808[0]));
  AL_DFF_0 al_d00399df (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21194118),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d72d808[1]));
  AL_DFF_0 al_d643feb4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2b6ee4f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d72d808[2]));
  AL_DFF_0 al_a71d5976 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fc2a0d6e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d72d808[3]));
  AL_DFF_0 al_cdc59d32 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_74d292d1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d72d808[4]));
  AL_DFF_0 al_9031820d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7ffa75b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d72d808[5]));
  AL_DFF_0 al_fce9ec32 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f76f90ba),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_905e5060[0]));
  AL_DFF_0 al_d2f60b9c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3cf942a1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_905e5060[1]));
  AL_DFF_0 al_87e7047d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e43903c1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_905e5060[2]));
  AL_DFF_0 al_c84ae31e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_512ab51),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_905e5060[3]));
  AL_DFF_0 al_40b79950 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3b1307c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_905e5060[4]));
  AL_DFF_0 al_e2201157 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b35f14e0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_905e5060[5]));
  AL_DFF_0 al_e66faf6a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4f5cc54),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62b22b32[0]));
  AL_DFF_0 al_931bcc2d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6a36379a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62b22b32[1]));
  AL_DFF_0 al_2fa9ec10 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_78cdcfba),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62b22b32[2]));
  AL_DFF_0 al_f096214d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_544aea7e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62b22b32[3]));
  AL_DFF_0 al_c291f35b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e9d913),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62b22b32[4]));
  AL_DFF_0 al_29a48406 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_20113785),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62b22b32[5]));
  AL_DFF_0 al_f276ec9e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_47c5e497),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f62f60e1[0]));
  AL_DFF_0 al_b4f3b6ab (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_42911267),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f62f60e1[1]));
  AL_DFF_0 al_6d7f2e4f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8abfdb0b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f62f60e1[2]));
  AL_DFF_0 al_e8a8c6dc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ce5ae5f4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f62f60e1[3]));
  AL_DFF_0 al_b76ed558 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3190947b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f62f60e1[4]));
  AL_DFF_0 al_85d61be8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a008bee3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f62f60e1[5]));
  AL_DFF_0 al_b981f636 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dce011d4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b737f75[0]));
  AL_DFF_0 al_174d41a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef04f6d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b737f75[1]));
  AL_DFF_0 al_8d42ca7d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71c5949d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b737f75[2]));
  AL_DFF_0 al_1ec50ee6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c721314),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b737f75[3]));
  AL_DFF_0 al_fc628718 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9cde5e3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b737f75[4]));
  AL_DFF_0 al_dd9d4c66 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_96bd601f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b737f75[5]));
  AL_DFF_0 al_3777b822 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b1f62da3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d7fecbad[0]));
  AL_DFF_0 al_2445bc4a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_42c99835),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d7fecbad[1]));
  AL_DFF_0 al_343f0014 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_800799cd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d7fecbad[2]));
  AL_DFF_0 al_3ffdc5e3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8f1d15d4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d7fecbad[3]));
  AL_DFF_0 al_30d7d295 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c6f34b3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d7fecbad[4]));
  AL_DFF_0 al_50f225b9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_85cc6a5c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d7fecbad[5]));
  AL_DFF_0 al_ea84d08d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2cb11ceb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d302088[0]));
  AL_DFF_0 al_ff9fa80f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bea784fd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d302088[1]));
  AL_DFF_0 al_efdc26b8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6b55c3b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d302088[2]));
  AL_DFF_0 al_db33796a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6169b199),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d302088[3]));
  AL_DFF_0 al_aaee18d5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d83b8ffa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d302088[4]));
  AL_DFF_0 al_c4f8ab1d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_26eb28a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d302088[5]));
  AL_DFF_0 al_81cba9f6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4ccae77b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_95e9fdd1[0]));
  AL_DFF_0 al_8feafca5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f33298c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_95e9fdd1[1]));
  AL_DFF_0 al_2afa3794 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b178800e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_95e9fdd1[2]));
  AL_DFF_0 al_39eabde7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef27da32),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_95e9fdd1[3]));
  AL_DFF_0 al_3dbe3b38 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ecb49f56),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_95e9fdd1[4]));
  AL_DFF_0 al_c83e135a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1eef59d6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_95e9fdd1[5]));
  AL_DFF_0 al_e9ba781a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_40c57b0a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_84027ae7[0]));
  AL_DFF_0 al_872b6e7d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f212ca88),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_84027ae7[1]));
  AL_DFF_0 al_c56228a9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7dedd4af),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_84027ae7[2]));
  AL_DFF_0 al_28aa7300 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_db2237d8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_84027ae7[3]));
  AL_DFF_0 al_fb373a9c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_688f86d6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_84027ae7[4]));
  AL_DFF_0 al_4bc32f62 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f9d8d0e0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_84027ae7[5]));
  AL_DFF_0 al_d818df07 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_59351be4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f61035a[0]));
  AL_DFF_0 al_6943780e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_697eb2f9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f61035a[1]));
  AL_DFF_0 al_e02ca4d6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_144891ce),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f61035a[2]));
  AL_DFF_0 al_28805c56 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c66c844),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f61035a[3]));
  AL_DFF_0 al_cf1f021a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d3983157),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f61035a[4]));
  AL_DFF_0 al_996ad3b9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_52ab1d02),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f61035a[5]));
  AL_DFF_0 al_1c5e946f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3fceb593),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4e28198f[0]));
  AL_DFF_0 al_95e2ce97 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2789af72),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4e28198f[1]));
  AL_DFF_0 al_869ebfaa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c803837c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4e28198f[2]));
  AL_DFF_0 al_ed1bb6c8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba93203f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4e28198f[3]));
  AL_DFF_0 al_d2dfb44 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1aca5917),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4e28198f[4]));
  AL_DFF_0 al_ce5fd90f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ca5bdee2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4e28198f[5]));
  AL_DFF_0 al_247b9835 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_806b722b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af419986[0]));
  AL_DFF_0 al_3f6585c0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d1caf9b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af419986[1]));
  AL_DFF_0 al_4e519c4a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_30f2f697),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af419986[2]));
  AL_DFF_0 al_43086caf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf317014),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af419986[3]));
  AL_DFF_0 al_7e1fe419 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_196ba081),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af419986[4]));
  AL_DFF_0 al_533683af (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba9d658c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af419986[5]));
  AL_DFF_0 al_ce9029ec (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3f65b31b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf0afe9a[0]));
  AL_DFF_0 al_89e5485e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_40a2a02d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf0afe9a[1]));
  AL_DFF_0 al_fe07d889 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_db637163),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf0afe9a[2]));
  AL_DFF_0 al_39e15326 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eaed5f24),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf0afe9a[3]));
  AL_DFF_0 al_2084fd1b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d82546f9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf0afe9a[4]));
  AL_DFF_0 al_bc5427ea (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_242f965e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf0afe9a[5]));
  AL_DFF_0 al_21d76be6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d0600950),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f594a8d9[0]));
  AL_DFF_0 al_65f3e37 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3ce57cf1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f594a8d9[1]));
  AL_DFF_0 al_f7b92890 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8d9fb1d7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f594a8d9[2]));
  AL_DFF_0 al_366ec005 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fc29ed6b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f594a8d9[3]));
  AL_DFF_0 al_43d8b97e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_61f6a76f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f594a8d9[4]));
  AL_DFF_0 al_8d03e341 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3b96714d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f594a8d9[5]));
  AL_DFF_0 al_ccb48ef6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f0955a51),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_df5cbc72[0]));
  AL_DFF_0 al_e2ed4aff (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3cbdf31),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_df5cbc72[1]));
  AL_DFF_0 al_63c2c1b9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4b874e94),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_df5cbc72[2]));
  AL_DFF_0 al_31451463 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_421da154),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_df5cbc72[3]));
  AL_DFF_0 al_58ac5e0e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_27924928),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_df5cbc72[4]));
  AL_DFF_0 al_56d7b6e5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_74987791),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_df5cbc72[5]));
  AL_DFF_0 al_89951133 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_855b52a9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdd95abd[0]));
  AL_DFF_0 al_47a71288 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_52e46bbb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdd95abd[1]));
  AL_DFF_0 al_4f167fc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8cc23669),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdd95abd[2]));
  AL_DFF_0 al_8dc29dd8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1e4cd67c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdd95abd[3]));
  AL_DFF_0 al_3310060c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d477830d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdd95abd[4]));
  AL_DFF_0 al_9d0c38b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff1bd228),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdd95abd[5]));
  AL_DFF_0 al_c05c2d4b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_353ab8af),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5d3b031[0]));
  AL_DFF_0 al_89a2cd65 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33e4a93b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5d3b031[1]));
  AL_DFF_0 al_af450579 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d4d15fe6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5d3b031[2]));
  AL_DFF_0 al_3e044440 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7bfa51e5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5d3b031[3]));
  AL_DFF_0 al_536db749 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ebef36bd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5d3b031[4]));
  AL_DFF_0 al_aefde2c6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f98cca52),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5d3b031[5]));
  AL_DFF_0 al_77e10335 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a5bb1940),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_79af3182[0]));
  AL_DFF_0 al_a9e50b10 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5bf1b92d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_79af3182[1]));
  AL_DFF_0 al_db7b9d69 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_14abcb2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_79af3182[2]));
  AL_DFF_0 al_474ee958 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_47108d32),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_79af3182[3]));
  AL_DFF_0 al_2b3deaca (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_91f0d008),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_79af3182[4]));
  AL_DFF_0 al_f29a63c2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dc467a61),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_79af3182[5]));
  AL_DFF_0 al_cbed9881 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5bce243b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_efab6074[0]));
  AL_DFF_0 al_aa82c2a2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_93118b48),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_efab6074[1]));
  AL_DFF_0 al_2836322b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef0d8a39),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_efab6074[2]));
  AL_DFF_0 al_14901cbb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_776135fb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_efab6074[3]));
  AL_DFF_0 al_6e3e8753 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fb7a2d43),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_efab6074[4]));
  AL_DFF_0 al_99099232 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c1ceb3d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_efab6074[5]));
  AL_DFF_0 al_42de6111 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2d7d45f8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6fdde80[0]));
  AL_DFF_0 al_ec1a5501 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_61210782),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6fdde80[1]));
  AL_DFF_0 al_4003d39e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c31bffdd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6fdde80[2]));
  AL_DFF_0 al_536f98a7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b265eaef),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6fdde80[3]));
  AL_DFF_0 al_50bd33f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2cea5c50),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6fdde80[4]));
  AL_DFF_0 al_3a366bc6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6263585f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6fdde80[5]));
  AL_DFF_0 al_c0b5827b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_efa11162),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e6b17901[0]));
  AL_DFF_0 al_b5ae2b8c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fe8d3a5b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e6b17901[1]));
  AL_DFF_0 al_7ac7a172 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_849ce6ee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e6b17901[2]));
  AL_DFF_0 al_fcf03899 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_67f1a13d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e6b17901[3]));
  AL_DFF_0 al_4320ed2d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef82c7c1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e6b17901[4]));
  AL_DFF_0 al_19641029 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_657419a5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e6b17901[5]));
  AL_DFF_0 al_50591232 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_462dcba0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57e2199e[0]));
  AL_DFF_0 al_c060308e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_13f4f154),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57e2199e[1]));
  AL_DFF_0 al_8962991d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1ec9bae4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57e2199e[2]));
  AL_DFF_0 al_a4d4ca17 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b87141aa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57e2199e[3]));
  AL_DFF_0 al_a9691a6a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7ebd1ee0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57e2199e[4]));
  AL_DFF_0 al_c67a117 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d735f43c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57e2199e[5]));
  AL_DFF_0 al_b98c07e7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d79f3cc5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48ac75ce[0]));
  AL_DFF_0 al_c494cc73 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_43d25c67),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48ac75ce[1]));
  AL_DFF_0 al_d863ce6d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4b9ffcd1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48ac75ce[2]));
  AL_DFF_0 al_48601094 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e690950c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48ac75ce[3]));
  AL_DFF_0 al_5b678efe (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55aa5549),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48ac75ce[4]));
  AL_DFF_0 al_63ff3f9d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_435a6ff0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48ac75ce[5]));
  AL_DFF_0 al_f2690062 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_24aa93c3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74387eee[0]));
  AL_DFF_0 al_5de4e9aa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4368302f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74387eee[1]));
  AL_DFF_0 al_667bb9fb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a9a47c58),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74387eee[2]));
  AL_DFF_0 al_9963d80c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bbf70a53),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74387eee[3]));
  AL_DFF_0 al_f1e30209 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_53cc11bb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74387eee[4]));
  AL_DFF_0 al_e55cb9bf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f7d22b96),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74387eee[5]));
  AL_DFF_0 al_c70c9f34 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7b6339b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7b20b0[0]));
  AL_DFF_0 al_9c127542 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d5903b66),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7b20b0[1]));
  AL_DFF_0 al_e5f2a457 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f9d6af3f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7b20b0[2]));
  AL_DFF_0 al_991e03f6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5d5a8704),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7b20b0[3]));
  AL_DFF_0 al_fb2d3e0a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b308bcff),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7b20b0[4]));
  AL_DFF_0 al_53d7f9bc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e14ba667),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7b20b0[5]));
  AL_DFF_0 al_3dade7e2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55e91735),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff281ad1[0]));
  AL_DFF_0 al_559efa81 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5edc286b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff281ad1[1]));
  AL_DFF_0 al_90f21c40 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_24cdfb7e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff281ad1[2]));
  AL_DFF_0 al_87b3e619 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_43e9197c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff281ad1[3]));
  AL_DFF_0 al_fb659afc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4966891e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff281ad1[4]));
  AL_DFF_0 al_7cf8526f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d196f7ed),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff281ad1[5]));
  AL_DFF_0 al_f390f42f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1b3ef09),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_effd30c4[0]));
  AL_DFF_0 al_3c59ddf2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3b949dc9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_effd30c4[1]));
  AL_DFF_0 al_d13f716a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3996c387),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_effd30c4[2]));
  AL_DFF_0 al_d53df85b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c792e14),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_effd30c4[3]));
  AL_DFF_0 al_eb31d198 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_40d3ac10),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_effd30c4[4]));
  AL_DFF_0 al_ad99c470 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e2d9e8f4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_effd30c4[5]));
  AL_DFF_0 al_d4fabc17 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_875e77a3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_adfe279[0]));
  AL_DFF_0 al_1299b7e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4afe32e3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_adfe279[1]));
  AL_DFF_0 al_aeaae454 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e841d4f6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_adfe279[2]));
  AL_DFF_0 al_2ef94d95 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7cd375ed),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_adfe279[3]));
  AL_DFF_0 al_cf8971ed (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e2b8e4f5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_adfe279[4]));
  AL_DFF_0 al_d4cf3bb7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fcebe00e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_adfe279[5]));
  AL_DFF_0 al_80c9e78f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dc060d66),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec6554e[0]));
  AL_DFF_0 al_fc27a3ec (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_37f1795f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec6554e[1]));
  AL_DFF_0 al_bfbe3ab0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6f9e8841),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec6554e[2]));
  AL_DFF_0 al_dcec5a34 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc31a928),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec6554e[3]));
  AL_DFF_0 al_39c0c1f7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3e845eb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec6554e[4]));
  AL_DFF_0 al_9d15f2b1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2be8e99),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec6554e[5]));
  AL_DFF_0 al_fe110a32 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e6bc3ac),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58c2706[0]));
  AL_DFF_0 al_af75acc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_59b8f11e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58c2706[1]));
  AL_DFF_0 al_19b918c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ca9ad4fa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58c2706[2]));
  AL_DFF_0 al_2b8a6fab (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b20e638),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58c2706[3]));
  AL_DFF_0 al_de4df651 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b39f3a2d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58c2706[4]));
  AL_DFF_0 al_87e75df9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2f8f631b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58c2706[5]));
  AL_DFF_0 al_95403baf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21e34e90),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1296b3[0]));
  AL_DFF_0 al_adb2406a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7e133bf5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1296b3[1]));
  AL_DFF_0 al_f5796ae8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ab7128ba),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1296b3[2]));
  AL_DFF_0 al_6da13b66 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_31b7b66),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1296b3[3]));
  AL_DFF_0 al_10d4a809 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_63dade5d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1296b3[4]));
  AL_DFF_0 al_ff56ac68 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a9bb616f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1296b3[5]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_6ec5044 (
    .a(al_31a603ae[0]),
    .b(al_527755ec[0]),
    .c(al_553ae5af[0]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_826c84b0));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_9681bbe7 (
    .a(al_826c84b0),
    .b(al_dd6ebfb0[0]),
    .c(al_81c227e0[0]),
    .o(al_5083706f));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_f373c0da (
    .a(al_31a603ae[3]),
    .b(al_527755ec[3]),
    .c(al_553ae5af[3]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_1c8bee0c));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_79f84c33 (
    .a(al_1c8bee0c),
    .b(al_dd6ebfb0[3]),
    .c(al_81c227e0[0]),
    .o(al_643bfe7d));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_db2df4c7 (
    .a(al_31a603ae[1]),
    .b(al_527755ec[1]),
    .c(al_553ae5af[1]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_12e98266));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_ca56921d (
    .a(al_12e98266),
    .b(al_dd6ebfb0[1]),
    .c(al_81c227e0[0]),
    .o(al_f6411514));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_94198fa0 (
    .a(al_31a603ae[2]),
    .b(al_527755ec[2]),
    .c(al_553ae5af[2]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_68fdf79b));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_a5056392 (
    .a(al_68fdf79b),
    .b(al_dd6ebfb0[2]),
    .c(al_81c227e0[0]),
    .o(al_6f628420));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*C*B*A)"),
    .INIT(64'h0000000080000000))
    al_7f2d3459 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_51a8d212));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*~D*~C*B*A)"),
    .INIT(64'h0000000000080000))
    al_dddef5f5 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_4706c253));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_34a4de84 (
    .a(al_31a603ae[4]),
    .b(al_527755ec[4]),
    .c(al_553ae5af[4]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_b05701c2));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_27795b5b (
    .a(al_b05701c2),
    .b(al_dd6ebfb0[4]),
    .c(al_81c227e0[0]),
    .o(al_95c3862c));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_83253e20 (
    .a(al_95c3862c),
    .b(al_4706c253),
    .c(al_84027ae7[4]),
    .o(al_688f86d6));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_f391b69 (
    .a(al_5083706f),
    .b(al_4706c253),
    .c(al_84027ae7[0]),
    .o(al_40c57b0a));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_5cbcf10a (
    .a(al_f6411514),
    .b(al_4706c253),
    .c(al_84027ae7[1]),
    .o(al_f212ca88));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_88a3fb32 (
    .a(al_6f628420),
    .b(al_4706c253),
    .c(al_84027ae7[2]),
    .o(al_7dedd4af));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_3da8ce3a (
    .a(al_643bfe7d),
    .b(al_4706c253),
    .c(al_84027ae7[3]),
    .o(al_db2237d8));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_f8d2171d (
    .a(al_4706c253),
    .b(al_84027ae7[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_f9d8d0e0));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*~C*B*A)"),
    .INIT(64'h0000000000000800))
    al_8134baaf (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_2e89ec2c));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_62ebb206 (
    .a(al_95c3862c),
    .b(al_2e89ec2c),
    .c(al_7b737f75[4]),
    .o(al_b9cde5e3));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_b639b3d7 (
    .a(al_5083706f),
    .b(al_2e89ec2c),
    .c(al_7b737f75[0]),
    .o(al_dce011d4));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e58fcc2b (
    .a(al_f6411514),
    .b(al_2e89ec2c),
    .c(al_7b737f75[1]),
    .o(al_ef04f6d));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1b9340c8 (
    .a(al_6f628420),
    .b(al_2e89ec2c),
    .c(al_7b737f75[2]),
    .o(al_71c5949d));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_72b74582 (
    .a(al_643bfe7d),
    .b(al_2e89ec2c),
    .c(al_7b737f75[3]),
    .o(al_c721314));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_1033b706 (
    .a(al_2e89ec2c),
    .b(al_7b737f75[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_96bd601f));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*~C*~B*A)"),
    .INIT(64'h0000020000000000))
    al_2c32748a (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_1d5f0c20));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1a1e71b3 (
    .a(al_95c3862c),
    .b(al_1d5f0c20),
    .c(al_a6fdde80[4]),
    .o(al_2cea5c50));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_f1a5e92 (
    .a(al_5083706f),
    .b(al_1d5f0c20),
    .c(al_a6fdde80[0]),
    .o(al_2d7d45f8));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_9f481eba (
    .a(al_f6411514),
    .b(al_1d5f0c20),
    .c(al_a6fdde80[1]),
    .o(al_61210782));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_b1568ea2 (
    .a(al_6f628420),
    .b(al_1d5f0c20),
    .c(al_a6fdde80[2]),
    .o(al_c31bffdd));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ae77f084 (
    .a(al_643bfe7d),
    .b(al_1d5f0c20),
    .c(al_a6fdde80[3]),
    .o(al_b265eaef));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_99683eb3 (
    .a(al_1d5f0c20),
    .b(al_a6fdde80[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_6263585f));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*~C*B*A)"),
    .INIT(64'h0800000000000000))
    al_ed086f56 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_a1fef711));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_55a64ee4 (
    .a(al_95c3862c),
    .b(al_a1fef711),
    .c(al_eec6554e[4]),
    .o(al_e3e845eb));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_18aed608 (
    .a(al_5083706f),
    .b(al_a1fef711),
    .c(al_eec6554e[0]),
    .o(al_dc060d66));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1e14b7e5 (
    .a(al_f6411514),
    .b(al_a1fef711),
    .c(al_eec6554e[1]),
    .o(al_37f1795f));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_350178ef (
    .a(al_6f628420),
    .b(al_a1fef711),
    .c(al_eec6554e[2]),
    .o(al_6f9e8841));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ad2a29e3 (
    .a(al_643bfe7d),
    .b(al_a1fef711),
    .c(al_eec6554e[3]),
    .o(al_bc31a928));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_1832126d (
    .a(al_a1fef711),
    .b(al_eec6554e[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_2be8e99));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_25953c2c (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_9ce674e2));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ae4dca09 (
    .a(al_95c3862c),
    .b(al_9ce674e2),
    .c(al_41bdf331[4]),
    .o(al_595cd185));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_571643c3 (
    .a(al_5083706f),
    .b(al_9ce674e2),
    .c(al_41bdf331[0]),
    .o(al_5b6e3903));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e3135a31 (
    .a(al_f6411514),
    .b(al_9ce674e2),
    .c(al_41bdf331[1]),
    .o(al_1f32b3ce));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_bbd9a9f3 (
    .a(al_6f628420),
    .b(al_9ce674e2),
    .c(al_41bdf331[2]),
    .o(al_4a3ec7d2));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_8fa73d80 (
    .a(al_643bfe7d),
    .b(al_9ce674e2),
    .c(al_41bdf331[3]),
    .o(al_1867b14e));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_2f859c86 (
    .a(al_9ce674e2),
    .b(al_41bdf331[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_d5c31119));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*~C*B*A)"),
    .INIT(64'h0000080000000000))
    al_50f7cc7 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_e7314734));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_9a8ecf65 (
    .a(al_95c3862c),
    .b(al_e7314734),
    .c(al_e6b17901[4]),
    .o(al_ef82c7c1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_d4263fe7 (
    .a(al_5083706f),
    .b(al_e7314734),
    .c(al_e6b17901[0]),
    .o(al_efa11162));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_cdef20f7 (
    .a(al_f6411514),
    .b(al_e7314734),
    .c(al_e6b17901[1]),
    .o(al_fe8d3a5b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_4df3a5f5 (
    .a(al_6f628420),
    .b(al_e7314734),
    .c(al_e6b17901[2]),
    .o(al_849ce6ee));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_418f6008 (
    .a(al_643bfe7d),
    .b(al_e7314734),
    .c(al_e6b17901[3]),
    .o(al_67f1a13d));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_2322b04e (
    .a(al_e7314734),
    .b(al_e6b17901[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_657419a5));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~D*C*~B*A)"),
    .INIT(64'h0020000000000000))
    al_33bf3e29 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_8ec42bd1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_cc0ebe40 (
    .a(al_95c3862c),
    .b(al_8ec42bd1),
    .c(al_ff281ad1[4]),
    .o(al_4966891e));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a87111ed (
    .a(al_5083706f),
    .b(al_8ec42bd1),
    .c(al_ff281ad1[0]),
    .o(al_55e91735));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_89e1de98 (
    .a(al_f6411514),
    .b(al_8ec42bd1),
    .c(al_ff281ad1[1]),
    .o(al_5edc286b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_3d95a827 (
    .a(al_6f628420),
    .b(al_8ec42bd1),
    .c(al_ff281ad1[2]),
    .o(al_24cdfb7e));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_43478be (
    .a(al_643bfe7d),
    .b(al_8ec42bd1),
    .c(al_ff281ad1[3]),
    .o(al_43e9197c));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_564a99db (
    .a(al_8ec42bd1),
    .b(al_ff281ad1[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_d196f7ed));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_1ec1536 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_754a5a85));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_fea7973 (
    .a(al_95c3862c),
    .b(al_754a5a85),
    .c(al_d7fecbad[4]),
    .o(al_c6f34b3));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_9700fdf8 (
    .a(al_5083706f),
    .b(al_754a5a85),
    .c(al_d7fecbad[0]),
    .o(al_b1f62da3));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_b43f8dff (
    .a(al_f6411514),
    .b(al_754a5a85),
    .c(al_d7fecbad[1]),
    .o(al_42c99835));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a7d04371 (
    .a(al_6f628420),
    .b(al_754a5a85),
    .c(al_d7fecbad[2]),
    .o(al_800799cd));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_c5bbe93c (
    .a(al_643bfe7d),
    .b(al_754a5a85),
    .c(al_d7fecbad[3]),
    .o(al_8f1d15d4));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_fa477db4 (
    .a(al_754a5a85),
    .b(al_d7fecbad[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_85cc6a5c));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*~B*A)"),
    .INIT(64'h2000000000000000))
    al_b739862d (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_86e6d7f8));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_b7960ca8 (
    .a(al_95c3862c),
    .b(al_86e6d7f8),
    .c(al_c58c2706[4]),
    .o(al_b39f3a2d));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_94639450 (
    .a(al_5083706f),
    .b(al_86e6d7f8),
    .c(al_c58c2706[0]),
    .o(al_3e6bc3ac));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a064129e (
    .a(al_f6411514),
    .b(al_86e6d7f8),
    .c(al_c58c2706[1]),
    .o(al_59b8f11e));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e4d57968 (
    .a(al_6f628420),
    .b(al_86e6d7f8),
    .c(al_c58c2706[2]),
    .o(al_ca9ad4fa));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_cf25abc5 (
    .a(al_643bfe7d),
    .b(al_86e6d7f8),
    .c(al_c58c2706[3]),
    .o(al_7b20e638));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_90c614ed (
    .a(al_86e6d7f8),
    .b(al_c58c2706[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_2f8f631b));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*~D*C*~B*A)"),
    .INIT(64'h0000000000200000))
    al_b45d5a2f (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_865f57bc));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_6da8bdea (
    .a(al_95c3862c),
    .b(al_865f57bc),
    .c(al_9f61035a[4]),
    .o(al_d3983157));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_4c850950 (
    .a(al_5083706f),
    .b(al_865f57bc),
    .c(al_9f61035a[0]),
    .o(al_59351be4));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_304b6751 (
    .a(al_f6411514),
    .b(al_865f57bc),
    .c(al_9f61035a[1]),
    .o(al_697eb2f9));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_2fbb7a05 (
    .a(al_6f628420),
    .b(al_865f57bc),
    .c(al_9f61035a[2]),
    .o(al_144891ce));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_fc65d885 (
    .a(al_643bfe7d),
    .b(al_865f57bc),
    .c(al_9f61035a[3]),
    .o(al_5c66c844));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_c18bd178 (
    .a(al_865f57bc),
    .b(al_9f61035a[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_52ab1d02));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_29bf4614 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_e54832a8));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_35cdea43 (
    .a(al_95c3862c),
    .b(al_e54832a8),
    .c(al_9d72d808[4]),
    .o(al_74d292d1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e524ceaa (
    .a(al_5083706f),
    .b(al_e54832a8),
    .c(al_9d72d808[0]),
    .o(al_dc426867));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_aae5743a (
    .a(al_f6411514),
    .b(al_e54832a8),
    .c(al_9d72d808[1]),
    .o(al_21194118));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_79403f56 (
    .a(al_6f628420),
    .b(al_e54832a8),
    .c(al_9d72d808[2]),
    .o(al_2b6ee4f));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_8c9497e0 (
    .a(al_643bfe7d),
    .b(al_e54832a8),
    .c(al_9d72d808[3]),
    .o(al_fc2a0d6e));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_f05d78d6 (
    .a(al_e54832a8),
    .b(al_9d72d808[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_7ffa75b1));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_3ea3b564 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_cd4f09bc));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_533443cc (
    .a(al_95c3862c),
    .b(al_cd4f09bc),
    .c(al_b1296b3[4]),
    .o(al_63dade5d));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_88bdb245 (
    .a(al_5083706f),
    .b(al_cd4f09bc),
    .c(al_b1296b3[0]),
    .o(al_21e34e90));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_226a2dc6 (
    .a(al_f6411514),
    .b(al_cd4f09bc),
    .c(al_b1296b3[1]),
    .o(al_7e133bf5));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_64202801 (
    .a(al_6f628420),
    .b(al_cd4f09bc),
    .c(al_b1296b3[2]),
    .o(al_ab7128ba));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_2f078df7 (
    .a(al_643bfe7d),
    .b(al_cd4f09bc),
    .c(al_b1296b3[3]),
    .o(al_31b7b66));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_bf248e81 (
    .a(al_cd4f09bc),
    .b(al_b1296b3[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_a9bb616f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*B*A)"),
    .INIT(64'h0000000000008000))
    al_e29a695b (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_a66b7d92));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_b4cd83b (
    .a(al_95c3862c),
    .b(al_a66b7d92),
    .c(al_8d302088[4]),
    .o(al_d83b8ffa));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a98fc2de (
    .a(al_5083706f),
    .b(al_a66b7d92),
    .c(al_8d302088[0]),
    .o(al_2cb11ceb));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_d8938aab (
    .a(al_f6411514),
    .b(al_a66b7d92),
    .c(al_8d302088[1]),
    .o(al_bea784fd));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_5d683fc0 (
    .a(al_6f628420),
    .b(al_a66b7d92),
    .c(al_8d302088[2]),
    .o(al_a6b55c3b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_7fef2e9a (
    .a(al_643bfe7d),
    .b(al_a66b7d92),
    .c(al_8d302088[3]),
    .o(al_6169b199));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_a93ffcfd (
    .a(al_a66b7d92),
    .b(al_8d302088[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_26eb28a));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*C*~B*A)"),
    .INIT(64'h0000002000000000))
    al_7a349979 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_364a5729));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_56999438 (
    .a(al_95c3862c),
    .b(al_364a5729),
    .c(al_79af3182[4]),
    .o(al_91f0d008));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_d5d1062 (
    .a(al_5083706f),
    .b(al_364a5729),
    .c(al_79af3182[0]),
    .o(al_a5bb1940));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_6f462c81 (
    .a(al_f6411514),
    .b(al_364a5729),
    .c(al_79af3182[1]),
    .o(al_5bf1b92d));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_5beb1c55 (
    .a(al_6f628420),
    .b(al_364a5729),
    .c(al_79af3182[2]),
    .o(al_14abcb2));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_84a135e3 (
    .a(al_643bfe7d),
    .b(al_364a5729),
    .c(al_79af3182[3]),
    .o(al_47108d32));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_f8232d5f (
    .a(al_364a5729),
    .b(al_79af3182[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_dc467a61));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*C*~B*A)"),
    .INIT(64'h0000000020000000))
    al_b423651f (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_fa88c9b1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1318aeae (
    .a(al_95c3862c),
    .b(al_fa88c9b1),
    .c(al_f594a8d9[4]),
    .o(al_61f6a76f));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_587400c7 (
    .a(al_5083706f),
    .b(al_fa88c9b1),
    .c(al_f594a8d9[0]),
    .o(al_d0600950));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ae033603 (
    .a(al_f6411514),
    .b(al_fa88c9b1),
    .c(al_f594a8d9[1]),
    .o(al_3ce57cf1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e1e2ded0 (
    .a(al_6f628420),
    .b(al_fa88c9b1),
    .c(al_f594a8d9[2]),
    .o(al_8d9fb1d7));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_328f6152 (
    .a(al_643bfe7d),
    .b(al_fa88c9b1),
    .c(al_f594a8d9[3]),
    .o(al_fc29ed6b));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_dd70dbf (
    .a(al_fa88c9b1),
    .b(al_f594a8d9[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_3b96714d));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*~D*C*B*A)"),
    .INIT(64'h0000000000800000))
    al_89f0c45e (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_d273ec64));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_77845e5 (
    .a(al_95c3862c),
    .b(al_d273ec64),
    .c(al_4e28198f[4]),
    .o(al_1aca5917));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_42fa719c (
    .a(al_5083706f),
    .b(al_d273ec64),
    .c(al_4e28198f[0]),
    .o(al_3fceb593));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_2ce6695a (
    .a(al_f6411514),
    .b(al_d273ec64),
    .c(al_4e28198f[1]),
    .o(al_2789af72));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e9e90801 (
    .a(al_6f628420),
    .b(al_d273ec64),
    .c(al_4e28198f[2]),
    .o(al_c803837c));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_6a8dba34 (
    .a(al_643bfe7d),
    .b(al_d273ec64),
    .c(al_4e28198f[3]),
    .o(al_ba93203f));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_f1b8f3f5 (
    .a(al_d273ec64),
    .b(al_4e28198f[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_ca5bdee2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*~B*A)"),
    .INIT(64'h0000000000000020))
    al_2d432e5d (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_29af3518));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ad7617a9 (
    .a(al_95c3862c),
    .b(al_29af3518),
    .c(al_905e5060[4]),
    .o(al_f3b1307c));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ada697a0 (
    .a(al_5083706f),
    .b(al_29af3518),
    .c(al_905e5060[0]),
    .o(al_f76f90ba));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a3ec16d1 (
    .a(al_f6411514),
    .b(al_29af3518),
    .c(al_905e5060[1]),
    .o(al_3cf942a1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1664289f (
    .a(al_6f628420),
    .b(al_29af3518),
    .c(al_905e5060[2]),
    .o(al_e43903c1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_312ba624 (
    .a(al_643bfe7d),
    .b(al_29af3518),
    .c(al_905e5060[3]),
    .o(al_512ab51));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_967c80a7 (
    .a(al_29af3518),
    .b(al_905e5060[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_b35f14e0));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*~D*~C*~B*A)"),
    .INIT(64'h0000000000020000))
    al_700fb4d8 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_27347df6));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a1621f56 (
    .a(al_95c3862c),
    .b(al_27347df6),
    .c(al_95e9fdd1[4]),
    .o(al_ecb49f56));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_8b4f270 (
    .a(al_5083706f),
    .b(al_27347df6),
    .c(al_95e9fdd1[0]),
    .o(al_4ccae77b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_687542ca (
    .a(al_f6411514),
    .b(al_27347df6),
    .c(al_95e9fdd1[1]),
    .o(al_f33298c));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ffaee60b (
    .a(al_6f628420),
    .b(al_27347df6),
    .c(al_95e9fdd1[2]),
    .o(al_b178800e));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_3133e58d (
    .a(al_643bfe7d),
    .b(al_27347df6),
    .c(al_95e9fdd1[3]),
    .o(al_ef27da32));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_94fe3096 (
    .a(al_27347df6),
    .b(al_95e9fdd1[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_1eef59d6));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*~C*~B*A)"),
    .INIT(64'h0200000000000000))
    al_fe29833d (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_b5aa848));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_c980a796 (
    .a(al_95c3862c),
    .b(al_b5aa848),
    .c(al_adfe279[4]),
    .o(al_e2b8e4f5));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_3d09dfca (
    .a(al_5083706f),
    .b(al_b5aa848),
    .c(al_adfe279[0]),
    .o(al_875e77a3));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_5f819a (
    .a(al_f6411514),
    .b(al_b5aa848),
    .c(al_adfe279[1]),
    .o(al_4afe32e3));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_f06bceb4 (
    .a(al_6f628420),
    .b(al_b5aa848),
    .c(al_adfe279[2]),
    .o(al_e841d4f6));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a55bb087 (
    .a(al_643bfe7d),
    .b(al_b5aa848),
    .c(al_adfe279[3]),
    .o(al_7cd375ed));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_af6ccf7f (
    .a(al_b5aa848),
    .b(al_adfe279[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_fcebe00e));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ac8ec86d (
    .a(al_95c3862c),
    .b(al_51a8d212),
    .c(al_df5cbc72[4]),
    .o(al_27924928));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1a3490f4 (
    .a(al_5083706f),
    .b(al_51a8d212),
    .c(al_df5cbc72[0]),
    .o(al_f0955a51));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_830416f3 (
    .a(al_f6411514),
    .b(al_51a8d212),
    .c(al_df5cbc72[1]),
    .o(al_c3cbdf31));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_828da705 (
    .a(al_6f628420),
    .b(al_51a8d212),
    .c(al_df5cbc72[2]),
    .o(al_4b874e94));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_920e2958 (
    .a(al_643bfe7d),
    .b(al_51a8d212),
    .c(al_df5cbc72[3]),
    .o(al_421da154));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_1f0235ba (
    .a(al_51a8d212),
    .b(al_df5cbc72[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_74987791));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~D*~C*~B*A)"),
    .INIT(64'h0002000000000000))
    al_6e3d63ef (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_1bfd1d5e));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_dbc06a82 (
    .a(al_95c3862c),
    .b(al_1bfd1d5e),
    .c(al_74387eee[4]),
    .o(al_53cc11bb));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_2741ebbb (
    .a(al_5083706f),
    .b(al_1bfd1d5e),
    .c(al_74387eee[0]),
    .o(al_24aa93c3));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_84c604ad (
    .a(al_f6411514),
    .b(al_1bfd1d5e),
    .c(al_74387eee[1]),
    .o(al_4368302f));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_6b31f335 (
    .a(al_6f628420),
    .b(al_1bfd1d5e),
    .c(al_74387eee[2]),
    .o(al_a9a47c58));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_83bdd76d (
    .a(al_643bfe7d),
    .b(al_1bfd1d5e),
    .c(al_74387eee[3]),
    .o(al_bbf70a53));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_23cce897 (
    .a(al_1bfd1d5e),
    .b(al_74387eee[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_f7d22b96));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*~C*~B*A)"),
    .INIT(64'h0000000002000000))
    al_f81ef50e (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_99e96d3e));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_d576e0cf (
    .a(al_95c3862c),
    .b(al_99e96d3e),
    .c(al_af419986[4]),
    .o(al_196ba081));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_771bd58c (
    .a(al_5083706f),
    .b(al_99e96d3e),
    .c(al_af419986[0]),
    .o(al_806b722b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_20a124c1 (
    .a(al_f6411514),
    .b(al_99e96d3e),
    .c(al_af419986[1]),
    .o(al_d1caf9b1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ddfdfadf (
    .a(al_6f628420),
    .b(al_99e96d3e),
    .c(al_af419986[2]),
    .o(al_30f2f697));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_bde152bb (
    .a(al_643bfe7d),
    .b(al_99e96d3e),
    .c(al_af419986[3]),
    .o(al_cf317014));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_c6a15cdc (
    .a(al_99e96d3e),
    .b(al_af419986[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_ba9d658c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*B*A)"),
    .INIT(64'h0000000000000080))
    al_122da31 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_5c28ad0a));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_f5ee80a (
    .a(al_95c3862c),
    .b(al_5c28ad0a),
    .c(al_62b22b32[4]),
    .o(al_e9d913));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ca1fbe8 (
    .a(al_5083706f),
    .b(al_5c28ad0a),
    .c(al_62b22b32[0]),
    .o(al_b4f5cc54));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a4f299e8 (
    .a(al_f6411514),
    .b(al_5c28ad0a),
    .c(al_62b22b32[1]),
    .o(al_6a36379a));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_63f713c1 (
    .a(al_6f628420),
    .b(al_5c28ad0a),
    .c(al_62b22b32[2]),
    .o(al_78cdcfba));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_156c5f9d (
    .a(al_643bfe7d),
    .b(al_5c28ad0a),
    .c(al_62b22b32[3]),
    .o(al_544aea7e));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_e6e0a15e (
    .a(al_5c28ad0a),
    .b(al_62b22b32[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_20113785));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~D*C*B*A)"),
    .INIT(64'h0080000000000000))
    al_57e3bbb4 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_fd33b43));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_17fe291c (
    .a(al_95c3862c),
    .b(al_fd33b43),
    .c(al_effd30c4[4]),
    .o(al_40d3ac10));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_3586dad5 (
    .a(al_5083706f),
    .b(al_fd33b43),
    .c(al_effd30c4[0]),
    .o(al_a1b3ef09));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ceeb9df5 (
    .a(al_f6411514),
    .b(al_fd33b43),
    .c(al_effd30c4[1]),
    .o(al_3b949dc9));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a60f8f54 (
    .a(al_6f628420),
    .b(al_fd33b43),
    .c(al_effd30c4[2]),
    .o(al_3996c387));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_8404223f (
    .a(al_643bfe7d),
    .b(al_fd33b43),
    .c(al_effd30c4[3]),
    .o(al_7c792e14));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_274894c1 (
    .a(al_fd33b43),
    .b(al_effd30c4[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_e2d9e8f4));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000200000000))
    al_67482e08 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_5c8dc62));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1280abbb (
    .a(al_95c3862c),
    .b(al_5c8dc62),
    .c(al_cdd95abd[4]),
    .o(al_d477830d));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_55e9d1ba (
    .a(al_5083706f),
    .b(al_5c8dc62),
    .c(al_cdd95abd[0]),
    .o(al_855b52a9));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_c3eaae1b (
    .a(al_f6411514),
    .b(al_5c8dc62),
    .c(al_cdd95abd[1]),
    .o(al_52e46bbb));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_2647b70b (
    .a(al_6f628420),
    .b(al_5c8dc62),
    .c(al_cdd95abd[2]),
    .o(al_8cc23669));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_feb046b4 (
    .a(al_643bfe7d),
    .b(al_5c8dc62),
    .c(al_cdd95abd[3]),
    .o(al_1e4cd67c));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_e86f026b (
    .a(al_5c8dc62),
    .b(al_cdd95abd[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_ff1bd228));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~D*~C*B*A)"),
    .INIT(64'h0008000000000000))
    al_1d53dfde (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_c1b01733));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_7bba0db0 (
    .a(al_95c3862c),
    .b(al_c1b01733),
    .c(al_c7b20b0[4]),
    .o(al_b308bcff));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_dcba48d7 (
    .a(al_5083706f),
    .b(al_c1b01733),
    .c(al_c7b20b0[0]),
    .o(al_b7b6339b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ea1e69fd (
    .a(al_f6411514),
    .b(al_c1b01733),
    .c(al_c7b20b0[1]),
    .o(al_d5903b66));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_9294e98f (
    .a(al_6f628420),
    .b(al_c1b01733),
    .c(al_c7b20b0[2]),
    .o(al_f9d6af3f));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_b06e075c (
    .a(al_643bfe7d),
    .b(al_c1b01733),
    .c(al_c7b20b0[3]),
    .o(al_5d5a8704));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_25d60317 (
    .a(al_c1b01733),
    .b(al_c7b20b0[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_e14ba667));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*C*B*A)"),
    .INIT(64'h0000800000000000))
    al_8f074ca3 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_dc901033));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_947d8a87 (
    .a(al_95c3862c),
    .b(al_dc901033),
    .c(al_48ac75ce[4]),
    .o(al_55aa5549));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1af57e1 (
    .a(al_5083706f),
    .b(al_dc901033),
    .c(al_48ac75ce[0]),
    .o(al_d79f3cc5));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_620ee42e (
    .a(al_f6411514),
    .b(al_dc901033),
    .c(al_48ac75ce[1]),
    .o(al_43d25c67));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_8a30c5ff (
    .a(al_6f628420),
    .b(al_dc901033),
    .c(al_48ac75ce[2]),
    .o(al_4b9ffcd1));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_dcd9317b (
    .a(al_643bfe7d),
    .b(al_dc901033),
    .c(al_48ac75ce[3]),
    .o(al_e690950c));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_d47f080e (
    .a(al_dc901033),
    .b(al_48ac75ce[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_435a6ff0));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*~C*B*A)"),
    .INIT(64'h0000000008000000))
    al_aac41bc5 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_53e4871));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_d5e3e06f (
    .a(al_95c3862c),
    .b(al_53e4871),
    .c(al_cf0afe9a[4]),
    .o(al_d82546f9));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_1009a8ab (
    .a(al_5083706f),
    .b(al_53e4871),
    .c(al_cf0afe9a[0]),
    .o(al_3f65b31b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_b37ee2c1 (
    .a(al_f6411514),
    .b(al_53e4871),
    .c(al_cf0afe9a[1]),
    .o(al_40a2a02d));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_af633b78 (
    .a(al_6f628420),
    .b(al_53e4871),
    .c(al_cf0afe9a[2]),
    .o(al_db637163));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_85387c1 (
    .a(al_643bfe7d),
    .b(al_53e4871),
    .c(al_cf0afe9a[3]),
    .o(al_eaed5f24));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_12e8a74d (
    .a(al_53e4871),
    .b(al_cf0afe9a[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_242f965e));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*~C*~B*A)"),
    .INIT(64'h0000000000000200))
    al_7d90ca46 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_5c9a1fe7));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e4c9c378 (
    .a(al_95c3862c),
    .b(al_5c9a1fe7),
    .c(al_f62f60e1[4]),
    .o(al_3190947b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_19f50554 (
    .a(al_5083706f),
    .b(al_5c9a1fe7),
    .c(al_f62f60e1[0]),
    .o(al_47c5e497));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_79492e92 (
    .a(al_f6411514),
    .b(al_5c9a1fe7),
    .c(al_f62f60e1[1]),
    .o(al_42911267));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_64e5ad87 (
    .a(al_6f628420),
    .b(al_5c9a1fe7),
    .c(al_f62f60e1[2]),
    .o(al_8abfdb0b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_cfce6dda (
    .a(al_643bfe7d),
    .b(al_5c9a1fe7),
    .c(al_f62f60e1[3]),
    .o(al_ce5ae5f4));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_816e12ba (
    .a(al_5c9a1fe7),
    .b(al_f62f60e1[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_a008bee3));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000800000000))
    al_543a54e0 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_317c528a));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e2a7c7dd (
    .a(al_95c3862c),
    .b(al_317c528a),
    .c(al_c5d3b031[4]),
    .o(al_ebef36bd));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_fd3ceb94 (
    .a(al_5083706f),
    .b(al_317c528a),
    .c(al_c5d3b031[0]),
    .o(al_353ab8af));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_8f11fef5 (
    .a(al_f6411514),
    .b(al_317c528a),
    .c(al_c5d3b031[1]),
    .o(al_33e4a93b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_18175678 (
    .a(al_6f628420),
    .b(al_317c528a),
    .c(al_c5d3b031[2]),
    .o(al_d4d15fe6));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ffff5a2d (
    .a(al_643bfe7d),
    .b(al_317c528a),
    .c(al_c5d3b031[3]),
    .o(al_7bfa51e5));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    al_dd8ca6af (
    .a(al_317c528a),
    .b(al_c5d3b031[5]),
    .c(al_81cbac46[0]),
    .d(al_81c227e0[0]),
    .o(al_f98cca52));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*C*B*A)"),
    .INIT(64'h0000008000000000))
    al_4b67d65 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_950c19d6));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_bccf4dc0 (
    .a(al_95c3862c),
    .b(al_950c19d6),
    .c(al_efab6074[4]),
    .o(al_fb7a2d43));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_613ae5e9 (
    .a(al_5083706f),
    .b(al_950c19d6),
    .c(al_efab6074[0]),
    .o(al_5bce243b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_82d4dee2 (
    .a(al_f6411514),
    .b(al_950c19d6),
    .c(al_efab6074[1]),
    .o(al_93118b48));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_e369134c (
    .a(al_6f628420),
    .b(al_950c19d6),
    .c(al_efab6074[2]),
    .o(al_ef0d8a39));
  AL_DFF_0 al_4f939a9d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_19acd84f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e1dd175[3]));
  AL_DFF_0 al_45e30107 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e097b175),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e1dd175[4]));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_3f207d2 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .f(al_5e1dd175[4]),
    .o(al_e097b175));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_d14da8d5 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .o(al_4b08729d));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    al_78ccdc26 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .o(al_153a7598));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*A))"),
    .INIT(16'h7f80))
    al_dda95744 (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .o(al_838dffd7));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*C*B*A))"),
    .INIT(32'h7fff8000))
    al_f81d3a0c (
    .a(al_9120ce24),
    .b(al_5e1dd175[0]),
    .c(al_5e1dd175[1]),
    .d(al_5e1dd175[2]),
    .e(al_5e1dd175[3]),
    .o(al_19acd84f));
  AL_DFF_0 al_4d3e8464 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4b08729d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e1dd175[0]));
  AL_DFF_0 al_4411c622 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_153a7598),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e1dd175[1]));
  AL_DFF_0 al_97e6e707 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_838dffd7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e1dd175[2]));
  AL_DFF_0 al_6a80b2be (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71c87c87[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_511af127[3]));
  AL_DFF_0 al_6fa25bf8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71c87c87[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_511af127[4]));
  AL_DFF_0 al_21309112 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71c87c87[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_511af127[0]));
  AL_DFF_0 al_f641777a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71c87c87[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_511af127[1]));
  AL_DFF_0 al_511393c5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71c87c87[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_511af127[2]));
  AL_DFF_0 al_a2c047cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[0]));
  AL_DFF_0 al_ef4904a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[1]));
  AL_DFF_0 al_ea6ba537 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[2]));
  AL_DFF_0 al_4d7cbb22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[3]));
  AL_DFF_0 al_e4842217 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[4]));
  AL_DFF_0 al_d41d97ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[5]));
  AL_DFF_0 al_36f8a011 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[6]));
  AL_DFF_0 al_87220067 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[7]));
  AL_DFF_0 al_ffcf5c9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[8]));
  AL_DFF_0 al_f6565c0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[9]));
  AL_DFF_0 al_583c5370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[10]));
  AL_DFF_0 al_664b2762 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[11]));
  AL_DFF_0 al_c463ac3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[12]));
  AL_DFF_0 al_ee9d20ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[13]));
  AL_DFF_0 al_c7707c82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[14]));
  AL_DFF_0 al_ec8414d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[15]));
  AL_DFF_0 al_da3ffce1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[16]));
  AL_DFF_0 al_377a86ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[17]));
  AL_DFF_0 al_9221265c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[18]));
  AL_DFF_0 al_67adf3dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[19]));
  AL_DFF_0 al_52c56d4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[20]));
  AL_DFF_0 al_bd6c2a7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[21]));
  AL_DFF_0 al_9e2e2ddf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[22]));
  AL_DFF_0 al_a70ee1ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[23]));
  AL_DFF_0 al_83fcf5be (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[24]));
  AL_DFF_0 al_c51991d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[25]));
  AL_DFF_0 al_aa9142dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[26]));
  AL_DFF_0 al_96640718 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[27]));
  AL_DFF_0 al_75ec1e71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[28]));
  AL_DFF_0 al_ad55bf83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[29]));
  AL_DFF_0 al_f1f6add6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[30]));
  AL_DFF_0 al_761c6697 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[31]));
  AL_DFF_0 al_7ca0fb57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[32]));
  AL_DFF_0 al_66a83c4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[33]));
  AL_DFF_0 al_6f33c0c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[34]));
  AL_DFF_0 al_d269dfd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[35]));
  AL_DFF_0 al_ae0d5461 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[36]));
  AL_DFF_0 al_f8866f8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[37]));
  AL_DFF_0 al_9e76cba2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[38]));
  AL_DFF_0 al_c386fb4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[39]));
  AL_DFF_0 al_5de2ee49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[40]));
  AL_DFF_0 al_8b4b2f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[41]));
  AL_DFF_0 al_164583c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[42]));
  AL_DFF_0 al_72b3c70c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[43]));
  AL_DFF_0 al_37b367f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[44]));
  AL_DFF_0 al_a7ca7c04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[45]));
  AL_DFF_0 al_83e1d787 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[46]));
  AL_DFF_0 al_121c3030 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[47]));
  AL_DFF_0 al_4bb44a4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[48]));
  AL_DFF_0 al_cb7456c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[49]));
  AL_DFF_0 al_f957bbad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[50]));
  AL_DFF_0 al_391d995e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[51]));
  AL_DFF_0 al_5da12c1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[52]));
  AL_DFF_0 al_69c04e37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[53]));
  AL_DFF_0 al_4b67da09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[54]));
  AL_DFF_0 al_d13d0c0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[55]));
  AL_DFF_0 al_336a790 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[56]));
  AL_DFF_0 al_4b92db75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[57]));
  AL_DFF_0 al_748b4493 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[58]));
  AL_DFF_0 al_7f8d5a15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[59]));
  AL_DFF_0 al_79771659 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[60]));
  AL_DFF_0 al_83ed60f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[61]));
  AL_DFF_0 al_2763b5cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[62]));
  AL_DFF_0 al_8f8634fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[63]));
  AL_DFF_0 al_c2bb7257 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[64]));
  AL_DFF_0 al_8573d509 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[65]));
  AL_DFF_0 al_b897a145 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[66]));
  AL_DFF_0 al_1f146f16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[67]));
  AL_DFF_0 al_2ea9c41c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[68]));
  AL_DFF_0 al_9a19c14a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[69]));
  AL_DFF_0 al_dfb38988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[70]));
  AL_DFF_0 al_526c6efb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[71]));
  AL_DFF_0 al_3778bf65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[72]));
  AL_DFF_0 al_c942afd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[73]));
  AL_DFF_0 al_3a68780 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[74]));
  AL_DFF_0 al_75deb3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[75]));
  AL_DFF_0 al_7b5c736e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[76]));
  AL_DFF_0 al_a98c1339 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[77]));
  AL_DFF_0 al_85f3e055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[78]));
  AL_DFF_0 al_f1b3b082 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[79]));
  AL_DFF_0 al_4eb96330 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[80]));
  AL_DFF_0 al_cfe9bcdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[81]));
  AL_DFF_0 al_f8745a53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[82]));
  AL_DFF_0 al_9306f5c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[83]));
  AL_DFF_0 al_7a65522a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[84]));
  AL_DFF_0 al_14d56ec7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[85]));
  AL_DFF_0 al_44c68a69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[86]));
  AL_DFF_0 al_5dc6b11d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[87]));
  AL_DFF_0 al_f81684fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[88]));
  AL_DFF_0 al_7e3e187d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[89]));
  AL_DFF_0 al_f9d2a488 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[90]));
  AL_DFF_0 al_94a2aa57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[91]));
  AL_DFF_0 al_fb382e77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[92]));
  AL_DFF_0 al_8530a059 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[93]));
  AL_DFF_0 al_35a4a392 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[94]));
  AL_DFF_0 al_e3494263 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[95]));
  AL_DFF_0 al_26063fef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[96]));
  AL_DFF_0 al_a590b464 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[97]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[97]));
  AL_DFF_0 al_6aa1ebb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[98]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[98]));
  AL_DFF_0 al_d5ff690 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[99]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[99]));
  AL_DFF_0 al_d3e5542b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[100]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[100]));
  AL_DFF_0 al_1fb5a5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[101]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[101]));
  AL_DFF_0 al_d5629505 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[102]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[102]));
  AL_DFF_0 al_d7ba2370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[103]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[103]));
  AL_DFF_0 al_e752d9b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[104]));
  AL_DFF_0 al_55776820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[105]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[105]));
  AL_DFF_0 al_a8385bcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[106]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[106]));
  AL_DFF_0 al_fe1743b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[107]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[107]));
  AL_DFF_0 al_7b838157 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[108]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[108]));
  AL_DFF_0 al_a0114bc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[109]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[109]));
  AL_DFF_0 al_9427f2a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[110]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[110]));
  AL_DFF_0 al_cb0352ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[111]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[111]));
  AL_DFF_0 al_767888fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[112]));
  AL_DFF_0 al_27ec2db1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[113]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[113]));
  AL_DFF_0 al_d7bdaed2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[114]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[114]));
  AL_DFF_0 al_526348ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[115]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[115]));
  AL_DFF_0 al_93ea114c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[116]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[116]));
  AL_DFF_0 al_abb12083 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[117]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[117]));
  AL_DFF_0 al_b0539ab2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[118]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[118]));
  AL_DFF_0 al_6293d1ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[119]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[119]));
  AL_DFF_0 al_94ebebbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[120]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[120]));
  AL_DFF_0 al_24b57da5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[121]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[121]));
  AL_DFF_0 al_61ea5f8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[122]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[122]));
  AL_DFF_0 al_40b40de5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[123]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[123]));
  AL_DFF_0 al_83300fa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[124]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[124]));
  AL_DFF_0 al_22a19530 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[125]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[125]));
  AL_DFF_0 al_7e372592 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[126]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[126]));
  AL_DFF_0 al_23095443 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[127]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[127]));
  AL_DFF_0 al_467676bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[128]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[128]));
  AL_DFF_0 al_19cf35e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[129]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[129]));
  AL_DFF_0 al_a13fae31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[130]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[130]));
  AL_DFF_0 al_1703c311 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[131]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[131]));
  AL_DFF_0 al_6b6918c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[132]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[132]));
  AL_DFF_0 al_445a9131 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[133]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[133]));
  AL_DFF_0 al_a46089c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[134]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[134]));
  AL_DFF_0 al_585bf2f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[135]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[135]));
  AL_DFF_0 al_6f64b202 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[136]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[136]));
  AL_DFF_0 al_611fbd76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[137]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[137]));
  AL_DFF_0 al_e9f3c556 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[138]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[138]));
  AL_DFF_0 al_7c61c41e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[139]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[139]));
  AL_DFF_0 al_7a97e545 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[140]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[140]));
  AL_DFF_0 al_b92fb102 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[141]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[141]));
  AL_DFF_0 al_e4c6a97a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[142]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[142]));
  AL_DFF_0 al_40520e6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[143]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[143]));
  AL_DFF_0 al_2ed8507b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[144]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[144]));
  AL_DFF_0 al_2b12a2a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[145]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[145]));
  AL_DFF_0 al_aebecaa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[146]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[146]));
  AL_DFF_0 al_eeb2779f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[147]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[147]));
  AL_DFF_0 al_b95176bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[148]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[148]));
  AL_DFF_0 al_28842731 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[149]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[149]));
  AL_DFF_0 al_d0a8147d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[150]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[150]));
  AL_DFF_0 al_f6dbecd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[151]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[151]));
  AL_DFF_0 al_5b62d487 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[152]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[152]));
  AL_DFF_0 al_f541018e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[153]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[153]));
  AL_DFF_0 al_e8b478f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[154]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[154]));
  AL_DFF_0 al_406a73f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[155]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[155]));
  AL_DFF_0 al_7fa31c69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[156]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[156]));
  AL_DFF_0 al_224f1266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[157]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[157]));
  AL_DFF_0 al_c9baa160 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[158]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[158]));
  AL_DFF_0 al_fa776952 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[159]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[159]));
  AL_DFF_0 al_52f8708c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[160]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[160]));
  AL_DFF_0 al_6fc5944 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[161]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[161]));
  AL_DFF_0 al_6c32e04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[162]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[162]));
  AL_DFF_0 al_5c63f54d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[163]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[163]));
  AL_DFF_0 al_415a738a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[164]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[164]));
  AL_DFF_0 al_645aad27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[165]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[165]));
  AL_DFF_0 al_4b7cc717 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[166]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[166]));
  AL_DFF_0 al_e4ae2b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[167]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[167]));
  AL_DFF_0 al_bc8bd9dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[168]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[168]));
  AL_DFF_0 al_f09493f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[169]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[169]));
  AL_DFF_0 al_21e3597e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[170]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[170]));
  AL_DFF_0 al_f9baccac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[171]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[171]));
  AL_DFF_0 al_54d5984c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[172]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[172]));
  AL_DFF_0 al_bcc87d2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[173]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[173]));
  AL_DFF_0 al_6d8fa2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[174]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[174]));
  AL_DFF_0 al_2f515552 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[175]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[175]));
  AL_DFF_0 al_b786be3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[176]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[176]));
  AL_DFF_0 al_78780ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[177]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[177]));
  AL_DFF_0 al_e8469c2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[178]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[178]));
  AL_DFF_0 al_29bd8365 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[179]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[179]));
  AL_DFF_0 al_e01d3465 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[180]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[180]));
  AL_DFF_0 al_e319446c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[181]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[181]));
  AL_DFF_0 al_a54b2fc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[182]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[182]));
  AL_DFF_0 al_605610f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[183]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[183]));
  AL_DFF_0 al_16cb5bc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[184]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[184]));
  AL_DFF_0 al_c15503f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[185]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[185]));
  AL_DFF_0 al_18dc9595 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[186]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[186]));
  AL_DFF_0 al_fe6b83b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[187]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[187]));
  AL_DFF_0 al_1f86e20e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[188]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[188]));
  AL_DFF_0 al_7a3edfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[189]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[189]));
  AL_DFF_0 al_707cc71f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[190]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[190]));
  AL_DFF_0 al_36575f50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[191]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[191]));
  AL_DFF_0 al_81cae855 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[192]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[192]));
  AL_DFF_0 al_4b15371f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[193]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[193]));
  AL_DFF_0 al_9b182cad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[194]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[194]));
  AL_DFF_0 al_297307bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[195]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[195]));
  AL_DFF_0 al_10fc63f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[196]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[196]));
  AL_DFF_0 al_15a28a86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[197]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[197]));
  AL_DFF_0 al_fe91b6d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[198]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[198]));
  AL_DFF_0 al_dbfc02ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[199]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[199]));
  AL_DFF_0 al_3adc9701 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[200]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[200]));
  AL_DFF_0 al_aa3636f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[201]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[201]));
  AL_DFF_0 al_c51e96f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[202]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[202]));
  AL_DFF_0 al_9114cd8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[203]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[203]));
  AL_DFF_0 al_9c83e0db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[204]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[204]));
  AL_DFF_0 al_98011877 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[205]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[205]));
  AL_DFF_0 al_302b55b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[206]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[206]));
  AL_DFF_0 al_ba7927dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[207]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[207]));
  AL_DFF_0 al_4ae60528 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[208]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[208]));
  AL_DFF_0 al_c211f239 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[209]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[209]));
  AL_DFF_0 al_f1702d8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[210]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[210]));
  AL_DFF_0 al_e2f78c36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[211]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[211]));
  AL_DFF_0 al_7ca0f11b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[212]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[212]));
  AL_DFF_0 al_89186bb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[213]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[213]));
  AL_DFF_0 al_1db9db30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[214]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[214]));
  AL_DFF_0 al_1833af60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[215]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[215]));
  AL_DFF_0 al_bd0ee853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[216]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[216]));
  AL_DFF_0 al_bd044e67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[217]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[217]));
  AL_DFF_0 al_b29058da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[218]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[218]));
  AL_DFF_0 al_9bf81fe8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[219]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[219]));
  AL_DFF_0 al_dd6094e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[220]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[220]));
  AL_DFF_0 al_9609e340 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[221]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[221]));
  AL_DFF_0 al_a025c545 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[222]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[222]));
  AL_DFF_0 al_214a0e16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[223]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[223]));
  AL_DFF_0 al_1fad7062 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[224]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[224]));
  AL_DFF_0 al_2b95c1b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[225]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[225]));
  AL_DFF_0 al_76ac6f28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[226]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[226]));
  AL_DFF_0 al_5beade04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[227]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[227]));
  AL_DFF_0 al_c94a7122 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[228]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[228]));
  AL_DFF_0 al_cd5ae007 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[229]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[229]));
  AL_DFF_0 al_c028056c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[230]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[230]));
  AL_DFF_0 al_1bbae4e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[231]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[231]));
  AL_DFF_0 al_a8bd263a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[232]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[232]));
  AL_DFF_0 al_a9fecaf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[233]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[233]));
  AL_DFF_0 al_49c39ae9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[234]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[234]));
  AL_DFF_0 al_17e1aee0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[235]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[235]));
  AL_DFF_0 al_b502a962 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[236]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[236]));
  AL_DFF_0 al_6aeff86f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[237]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[237]));
  AL_DFF_0 al_1476349d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[238]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[238]));
  AL_DFF_0 al_a7363e8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[239]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[239]));
  AL_DFF_0 al_9504ec73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[240]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[240]));
  AL_DFF_0 al_3f0133a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[241]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[241]));
  AL_DFF_0 al_a69a700c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[242]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[242]));
  AL_DFF_0 al_64955697 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[243]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[243]));
  AL_DFF_0 al_e3f66dc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[244]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[244]));
  AL_DFF_0 al_bc52eaf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[245]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[245]));
  AL_DFF_0 al_5e2a9bc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[246]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[246]));
  AL_DFF_0 al_20cfb3d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[247]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[247]));
  AL_DFF_0 al_2dcbcde7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[248]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[248]));
  AL_DFF_0 al_840d6c96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[249]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[249]));
  AL_DFF_0 al_17a7a44f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[250]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[250]));
  AL_DFF_0 al_a11bade7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[251]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[251]));
  AL_DFF_0 al_cf30af9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[252]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[252]));
  AL_DFF_0 al_d16ad1fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[253]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[253]));
  AL_DFF_0 al_15896eb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[254]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[254]));
  AL_DFF_0 al_70365442 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1952ddef[255]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31a3e7af[255]));
  AL_DFF_0 al_6b253a30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[0]));
  AL_DFF_0 al_20a419da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[1]));
  AL_DFF_0 al_765ab5fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[2]));
  AL_DFF_0 al_9fbb3345 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[3]));
  AL_DFF_0 al_3a416326 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[4]));
  AL_DFF_0 al_9d0789a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[5]));
  AL_DFF_0 al_6479ae4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[6]));
  AL_DFF_0 al_f69f5c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[7]));
  AL_DFF_0 al_8e5ec9d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[8]));
  AL_DFF_0 al_a388dd00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[9]));
  AL_DFF_0 al_fb46f3f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[10]));
  AL_DFF_0 al_eb24d16d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[11]));
  AL_DFF_0 al_609c1200 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[12]));
  AL_DFF_0 al_fdf3f6a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[13]));
  AL_DFF_0 al_47b28d59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[14]));
  AL_DFF_0 al_4b323199 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[15]));
  AL_DFF_0 al_d65c07c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[16]));
  AL_DFF_0 al_9f3a008e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[17]));
  AL_DFF_0 al_cd7048f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[18]));
  AL_DFF_0 al_32a14a4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[19]));
  AL_DFF_0 al_177d6710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[20]));
  AL_DFF_0 al_380191d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[21]));
  AL_DFF_0 al_8a83705a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[22]));
  AL_DFF_0 al_ea1edb89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[23]));
  AL_DFF_0 al_988ba4be (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[24]));
  AL_DFF_0 al_bfb3386b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[97]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[25]));
  AL_DFF_0 al_458b8fbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[98]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[26]));
  AL_DFF_0 al_d6b68f44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[99]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[27]));
  AL_DFF_0 al_a5ed1724 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[100]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[28]));
  AL_DFF_0 al_14226e96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[101]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[29]));
  AL_DFF_0 al_3a51ac47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[102]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[30]));
  AL_DFF_0 al_f1b500d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[103]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[31]));
  AL_DFF_0 al_a0731037 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[128]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[32]));
  AL_DFF_0 al_71ca5882 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[129]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[33]));
  AL_DFF_0 al_ff6425ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[130]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[34]));
  AL_DFF_0 al_30ec1327 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[131]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[35]));
  AL_DFF_0 al_352bc939 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[132]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[36]));
  AL_DFF_0 al_7e4d597f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[133]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[37]));
  AL_DFF_0 al_771aaf75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[134]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[38]));
  AL_DFF_0 al_3b03124b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[135]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[39]));
  AL_DFF_0 al_7b87c997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[160]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[40]));
  AL_DFF_0 al_5b564dd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[161]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[41]));
  AL_DFF_0 al_86e5f36d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[162]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[42]));
  AL_DFF_0 al_46ff90d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[163]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[43]));
  AL_DFF_0 al_a030329a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[164]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[44]));
  AL_DFF_0 al_f6b7f7b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[165]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[45]));
  AL_DFF_0 al_82de6767 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[166]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[46]));
  AL_DFF_0 al_2c02f355 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[167]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[47]));
  AL_DFF_0 al_4e1fdcab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[192]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[48]));
  AL_DFF_0 al_fc3a179e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[193]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[49]));
  AL_DFF_0 al_8a11a27e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[194]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[50]));
  AL_DFF_0 al_c09e10a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[195]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[51]));
  AL_DFF_0 al_e507bc75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[196]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[52]));
  AL_DFF_0 al_2d8ad5e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[197]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[53]));
  AL_DFF_0 al_3fd20942 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[198]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[54]));
  AL_DFF_0 al_2458f70d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[199]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[55]));
  AL_DFF_0 al_612a46e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[224]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[56]));
  AL_DFF_0 al_642b0cc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[225]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[57]));
  AL_DFF_0 al_a63426a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[226]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[58]));
  AL_DFF_0 al_ab525067 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[227]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[59]));
  AL_DFF_0 al_b0b17bf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[228]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[60]));
  AL_DFF_0 al_63407262 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[229]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[61]));
  AL_DFF_0 al_edba2cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[230]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[62]));
  AL_DFF_0 al_d6ac2f1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[231]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[63]));
  AL_DFF_0 al_c31f927b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[64]));
  AL_DFF_0 al_cbbf1ae6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[65]));
  AL_DFF_0 al_3ddb928a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[66]));
  AL_DFF_0 al_cc49a379 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[67]));
  AL_DFF_0 al_40371286 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[68]));
  AL_DFF_0 al_130d6542 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[69]));
  AL_DFF_0 al_40ab55c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[70]));
  AL_DFF_0 al_54322eb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[71]));
  AL_DFF_0 al_7c9e6fe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[72]));
  AL_DFF_0 al_aa211768 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[73]));
  AL_DFF_0 al_ff8be249 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[74]));
  AL_DFF_0 al_37107d91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[75]));
  AL_DFF_0 al_31c6c01a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[76]));
  AL_DFF_0 al_36d24647 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[77]));
  AL_DFF_0 al_ed9cec90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[78]));
  AL_DFF_0 al_b80d1593 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[79]));
  AL_DFF_0 al_f322783c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[80]));
  AL_DFF_0 al_701f46ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[81]));
  AL_DFF_0 al_c2c77052 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[82]));
  AL_DFF_0 al_7a8d2728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[83]));
  AL_DFF_0 al_b09bc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[84]));
  AL_DFF_0 al_364d3371 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[85]));
  AL_DFF_0 al_9a7ebdad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[86]));
  AL_DFF_0 al_2237591e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[87]));
  AL_DFF_0 al_2e69b7c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[88]));
  AL_DFF_0 al_ff7020f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[105]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[89]));
  AL_DFF_0 al_281c01bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[106]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[90]));
  AL_DFF_0 al_ff386a17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[107]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[91]));
  AL_DFF_0 al_738755ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[108]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[92]));
  AL_DFF_0 al_a016b5cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[109]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[93]));
  AL_DFF_0 al_26b94a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[110]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[94]));
  AL_DFF_0 al_50d73bcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[111]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[95]));
  AL_DFF_0 al_4909f420 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[136]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[96]));
  AL_DFF_0 al_5cf0b3e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[137]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[97]));
  AL_DFF_0 al_fb2d7256 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[138]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[98]));
  AL_DFF_0 al_ee84d6e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[139]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[99]));
  AL_DFF_0 al_5b43e8cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[140]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[100]));
  AL_DFF_0 al_e7b1a4f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[141]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[101]));
  AL_DFF_0 al_d51fcc96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[142]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[102]));
  AL_DFF_0 al_782a4c79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[143]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[103]));
  AL_DFF_0 al_fd3ae05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[168]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[104]));
  AL_DFF_0 al_4d1e45be (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[169]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[105]));
  AL_DFF_0 al_c384d4cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[170]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[106]));
  AL_DFF_0 al_95bab56c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[171]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[107]));
  AL_DFF_0 al_e0c05aa3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[172]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[108]));
  AL_DFF_0 al_67b933ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[173]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[109]));
  AL_DFF_0 al_b0bf6cff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[174]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[110]));
  AL_DFF_0 al_bebd1e1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[175]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[111]));
  AL_DFF_0 al_2f428a7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[200]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[112]));
  AL_DFF_0 al_c39726c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[201]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[113]));
  AL_DFF_0 al_20d512e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[202]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[114]));
  AL_DFF_0 al_fa7e1fa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[203]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[115]));
  AL_DFF_0 al_dcdff0a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[204]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[116]));
  AL_DFF_0 al_63cbc825 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[205]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[117]));
  AL_DFF_0 al_cacb16e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[206]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[118]));
  AL_DFF_0 al_b7f865e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[207]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[119]));
  AL_DFF_0 al_4a7cf84b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[232]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[120]));
  AL_DFF_0 al_b90d2e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[233]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[121]));
  AL_DFF_0 al_d5472126 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[234]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[122]));
  AL_DFF_0 al_276ce216 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[235]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[123]));
  AL_DFF_0 al_f2e3d69a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[236]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[124]));
  AL_DFF_0 al_fd330492 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[237]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[125]));
  AL_DFF_0 al_69eda7e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[238]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[126]));
  AL_DFF_0 al_844b4486 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[239]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[127]));
  AL_DFF_0 al_137d7592 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[128]));
  AL_DFF_0 al_c92263ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[129]));
  AL_DFF_0 al_b34e970a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[130]));
  AL_DFF_0 al_c9274bcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[131]));
  AL_DFF_0 al_bb013c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[132]));
  AL_DFF_0 al_1932cd5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[133]));
  AL_DFF_0 al_19d01433 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[134]));
  AL_DFF_0 al_2a2eb0ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[135]));
  AL_DFF_0 al_44be74bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[136]));
  AL_DFF_0 al_6c529ea9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[137]));
  AL_DFF_0 al_5049017d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[138]));
  AL_DFF_0 al_e9101607 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[139]));
  AL_DFF_0 al_f287cf51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[140]));
  AL_DFF_0 al_affdb86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[141]));
  AL_DFF_0 al_ee114b04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[142]));
  AL_DFF_0 al_9633677d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[143]));
  AL_DFF_0 al_2d9aa43c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[144]));
  AL_DFF_0 al_a2ada479 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[145]));
  AL_DFF_0 al_e1fbf09c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[146]));
  AL_DFF_0 al_821c15d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[147]));
  AL_DFF_0 al_17d6bab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[148]));
  AL_DFF_0 al_c0f69cac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[149]));
  AL_DFF_0 al_6a439cb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[150]));
  AL_DFF_0 al_a5e49158 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[151]));
  AL_DFF_0 al_43f214da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[152]));
  AL_DFF_0 al_6745f674 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[113]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[153]));
  AL_DFF_0 al_d5ba7c40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[114]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[154]));
  AL_DFF_0 al_ae0a723d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[115]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[155]));
  AL_DFF_0 al_430e4215 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[116]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[156]));
  AL_DFF_0 al_ca3e1f36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[117]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[157]));
  AL_DFF_0 al_a66856ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[118]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[158]));
  AL_DFF_0 al_21bd9f3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[119]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[159]));
  AL_DFF_0 al_202d6a5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[144]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[160]));
  AL_DFF_0 al_66919bef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[145]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[161]));
  AL_DFF_0 al_2275d0c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[146]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[162]));
  AL_DFF_0 al_35950dff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[147]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[163]));
  AL_DFF_0 al_f12b10a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[148]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[164]));
  AL_DFF_0 al_66b9e50b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[149]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[165]));
  AL_DFF_0 al_ffb93dc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[150]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[166]));
  AL_DFF_0 al_2b0ba2f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[151]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[167]));
  AL_DFF_0 al_db34dd31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[176]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[168]));
  AL_DFF_0 al_77ae4e02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[177]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[169]));
  AL_DFF_0 al_8b145ead (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[178]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[170]));
  AL_DFF_0 al_bebe7e38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[179]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[171]));
  AL_DFF_0 al_cb098cce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[180]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[172]));
  AL_DFF_0 al_9931c301 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[181]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[173]));
  AL_DFF_0 al_32f8085b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[182]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[174]));
  AL_DFF_0 al_d94c8b2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[183]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[175]));
  AL_DFF_0 al_17902b63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[208]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[176]));
  AL_DFF_0 al_52f9e320 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[209]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[177]));
  AL_DFF_0 al_f2e9aa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[210]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[178]));
  AL_DFF_0 al_88a333e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[211]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[179]));
  AL_DFF_0 al_89d568cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[212]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[180]));
  AL_DFF_0 al_7cf88b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[213]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[181]));
  AL_DFF_0 al_8a512fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[214]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[182]));
  AL_DFF_0 al_874bc148 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[215]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[183]));
  AL_DFF_0 al_9b5e468b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[240]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[184]));
  AL_DFF_0 al_77e7eb92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[241]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[185]));
  AL_DFF_0 al_ac789c3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[242]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[186]));
  AL_DFF_0 al_80d5d359 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[243]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[187]));
  AL_DFF_0 al_834b5f9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[244]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[188]));
  AL_DFF_0 al_be4dcd0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[245]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[189]));
  AL_DFF_0 al_89e8ea24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[246]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[190]));
  AL_DFF_0 al_aabcdc38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[247]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[191]));
  AL_DFF_0 al_4cb33297 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[192]));
  AL_DFF_0 al_dda4de4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[193]));
  AL_DFF_0 al_8a45f99d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[194]));
  AL_DFF_0 al_a992caa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[195]));
  AL_DFF_0 al_aa7efa28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[196]));
  AL_DFF_0 al_1f1009eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[197]));
  AL_DFF_0 al_28619e99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[198]));
  AL_DFF_0 al_bd40f0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[199]));
  AL_DFF_0 al_c6895aaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[200]));
  AL_DFF_0 al_2618698f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[201]));
  AL_DFF_0 al_6c68791b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[202]));
  AL_DFF_0 al_c1cc5a13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[203]));
  AL_DFF_0 al_61cfc573 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[204]));
  AL_DFF_0 al_c41ccdce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[205]));
  AL_DFF_0 al_c60cab6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[206]));
  AL_DFF_0 al_c0b684b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[207]));
  AL_DFF_0 al_31865243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[208]));
  AL_DFF_0 al_a2362c6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[209]));
  AL_DFF_0 al_b854cb0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[210]));
  AL_DFF_0 al_2c0d953 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[211]));
  AL_DFF_0 al_44615df8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[212]));
  AL_DFF_0 al_11ca59ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[213]));
  AL_DFF_0 al_b4cbd241 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[214]));
  AL_DFF_0 al_2d1a64b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[215]));
  AL_DFF_0 al_63c7ce58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[120]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[216]));
  AL_DFF_0 al_401ede44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[121]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[217]));
  AL_DFF_0 al_ee1bf9da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[122]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[218]));
  AL_DFF_0 al_ba990dbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[123]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[219]));
  AL_DFF_0 al_2af6dab0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[124]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[220]));
  AL_DFF_0 al_16119147 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[125]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[221]));
  AL_DFF_0 al_1f0a1243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[126]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[222]));
  AL_DFF_0 al_16e68506 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[127]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[223]));
  AL_DFF_0 al_8d743085 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[152]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[224]));
  AL_DFF_0 al_d7f2f1c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[153]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[225]));
  AL_DFF_0 al_cfce363a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[154]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[226]));
  AL_DFF_0 al_2cfed5c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[155]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[227]));
  AL_DFF_0 al_7219a51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[156]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[228]));
  AL_DFF_0 al_6613fb66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[157]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[229]));
  AL_DFF_0 al_b28dfa61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[158]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[230]));
  AL_DFF_0 al_658b6c5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[159]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[231]));
  AL_DFF_0 al_ef241f99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[184]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[232]));
  AL_DFF_0 al_fca4571b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[185]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[233]));
  AL_DFF_0 al_7ab1bcf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[186]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[234]));
  AL_DFF_0 al_4a2a4901 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[187]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[235]));
  AL_DFF_0 al_adecc544 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[188]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[236]));
  AL_DFF_0 al_5bc45b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[189]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[237]));
  AL_DFF_0 al_ad785af5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[190]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[238]));
  AL_DFF_0 al_9d1addc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[191]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[239]));
  AL_DFF_0 al_4e72bd8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[216]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[240]));
  AL_DFF_0 al_92713a31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[217]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[241]));
  AL_DFF_0 al_6fef3347 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[218]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[242]));
  AL_DFF_0 al_eaff99a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[219]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[243]));
  AL_DFF_0 al_8d9aca9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[220]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[244]));
  AL_DFF_0 al_740bf220 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[221]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[245]));
  AL_DFF_0 al_762595b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[222]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[246]));
  AL_DFF_0 al_15e94601 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[223]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[247]));
  AL_DFF_0 al_6dee98ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[248]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[248]));
  AL_DFF_0 al_d6d2925d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[249]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[249]));
  AL_DFF_0 al_f61f7b2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[250]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[250]));
  AL_DFF_0 al_54894f74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[251]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[251]));
  AL_DFF_0 al_2f9573b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[252]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[252]));
  AL_DFF_0 al_70f6b7ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[253]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[253]));
  AL_DFF_0 al_fb292df4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[254]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[254]));
  AL_DFF_0 al_17d6cc11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(dfi_rddata_w[255]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1952ddef[255]));
  AL_DFF_0 al_914fc3ca (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0f3a3cd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0f3a3cd[0]));
  AL_DFF_0 al_441d6163 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0f3a3cd[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0f3a3cd[2]));
  AL_DFF_0 al_71e5e181 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4aabc590[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0f3a3cd[3]));
  AL_DFF_0 al_879f22cb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4aabc590[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0f3a3cd[6]));
  AL_DFF_0 al_b508d810 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4aabc590[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0f3a3cd[7]));
  AL_DFF_0 al_87337529 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_83bf73ec),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af133298[0]));
  AL_DFF_0 al_d42994de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_342187f3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af133298[1]));
  AL_DFF_0 al_1f40eef4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4cf135b8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af133298[2]));
  AL_DFF_0 al_e3da6788 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9aab1a4f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af133298[3]));
  AL_DFF_0 al_a22b15ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_af133298[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af133298[5]));
  AL_DFF_0 al_8a28b6a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_af133298[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af133298[6]));
  AL_DFF_0 al_15704778 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_af133298[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af133298[7]));
  AL_DFF_0 al_25fb7e75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_af133298[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af133298[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d1cbea55 (
    .a(al_5083706f),
    .b(al_ef9accde),
    .o(al_83bf73ec));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_8efca354 (
    .a(al_643bfe7d),
    .b(al_ef9accde),
    .o(al_9aab1a4f));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_607272fa (
    .a(al_f6411514),
    .b(al_ef9accde),
    .o(al_342187f3));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_42515022 (
    .a(al_6f628420),
    .b(al_ef9accde),
    .o(al_4cf135b8));
  AL_DFF_0 al_fab3677 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[0]));
  AL_DFF_0 al_73c24240 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[1]));
  AL_DFF_0 al_9a5a345 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[2]));
  AL_DFF_0 al_f4cdba6c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[3]));
  AL_DFF_0 al_c7ca4f2b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[4]));
  AL_DFF_0 al_b4f84c14 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[5]));
  AL_DFF_0 al_8b4afbc2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[6]));
  AL_DFF_0 al_aa8330ad (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[7]));
  AL_DFF_0 al_63d48c70 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[32]));
  AL_DFF_0 al_1bede9f1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[33]));
  AL_DFF_0 al_489b4618 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[34]));
  AL_DFF_0 al_a6fece49 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[35]));
  AL_DFF_0 al_74171de8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[36]));
  AL_DFF_0 al_3eb73f5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[37]));
  AL_DFF_0 al_ed14c142 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[38]));
  AL_DFF_0 al_f8baf227 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[39]));
  AL_DFF_0 al_9440f517 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[64]));
  AL_DFF_0 al_8487ecb3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[65]));
  AL_DFF_0 al_906843bb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[66]));
  AL_DFF_0 al_c7b936dc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[67]));
  AL_DFF_0 al_85c7c358 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[68]));
  AL_DFF_0 al_3afc29d1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[69]));
  AL_DFF_0 al_7176e400 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[70]));
  AL_DFF_0 al_a29aa681 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[71]));
  AL_DFF_0 al_c18ada98 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[96]));
  AL_DFF_0 al_ab27fc39 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[97]));
  AL_DFF_0 al_5279d7a3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[98]));
  AL_DFF_0 al_56500611 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[99]));
  AL_DFF_0 al_94852772 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[100]));
  AL_DFF_0 al_417a8bb7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[101]));
  AL_DFF_0 al_7c9d04a5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[102]));
  AL_DFF_0 al_fee1ba20 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32e78cf2[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[103]));
  AL_DFF_0 al_5f58593a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[128]));
  AL_DFF_0 al_5276553a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[129]));
  AL_DFF_0 al_eee73b64 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[130]));
  AL_DFF_0 al_4ca045bc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[131]));
  AL_DFF_0 al_8e1d287d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[132]));
  AL_DFF_0 al_791dc526 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[133]));
  AL_DFF_0 al_33dc8061 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[134]));
  AL_DFF_0 al_c805fd69 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[135]));
  AL_DFF_0 al_6b2f3d7d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[160]));
  AL_DFF_0 al_eed8037 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[161]));
  AL_DFF_0 al_d76cadc5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[162]));
  AL_DFF_0 al_73124b56 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[163]));
  AL_DFF_0 al_b660030d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[164]));
  AL_DFF_0 al_dff6d388 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[165]));
  AL_DFF_0 al_96b16488 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[166]));
  AL_DFF_0 al_2ae31a78 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[167]));
  AL_DFF_0 al_bbf51030 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[192]));
  AL_DFF_0 al_9e3d5f02 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[193]));
  AL_DFF_0 al_276f58a5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[194]));
  AL_DFF_0 al_ba490cb7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[195]));
  AL_DFF_0 al_6c31368d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[196]));
  AL_DFF_0 al_1f90af31 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[197]));
  AL_DFF_0 al_1435e63d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[198]));
  AL_DFF_0 al_7c490b1f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[199]));
  AL_DFF_0 al_a169c888 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[224]));
  AL_DFF_0 al_b3653cc5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[225]));
  AL_DFF_0 al_ba0fc02c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[226]));
  AL_DFF_0 al_2f2e1481 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[227]));
  AL_DFF_0 al_28de05f9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[228]));
  AL_DFF_0 al_b84a3bda (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[229]));
  AL_DFF_0 al_c1e21d4e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[230]));
  AL_DFF_0 al_c327a0c1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[231]));
  AL_DFF_0 al_a8e69747 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[64]));
  AL_DFF_0 al_40c82c97 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[65]));
  AL_DFF_0 al_ea402be7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[66]));
  AL_DFF_0 al_68ae6d33 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[67]));
  AL_DFF_0 al_257e6483 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[68]));
  AL_DFF_0 al_3ff4a082 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[69]));
  AL_DFF_0 al_61260ff0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[70]));
  AL_DFF_0 al_ee8e150e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[71]));
  AL_DFF_0 al_f2b17265 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[72]));
  AL_DFF_0 al_202f4e10 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[73]));
  AL_DFF_0 al_f8f76c1b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[74]));
  AL_DFF_0 al_707ba85a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[75]));
  AL_DFF_0 al_b2ccf1f2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[76]));
  AL_DFF_0 al_37d884a9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[77]));
  AL_DFF_0 al_5aa05ad3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[78]));
  AL_DFF_0 al_8f3e9484 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[79]));
  AL_DFF_0 al_880ff29b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[80]));
  AL_DFF_0 al_8afca97 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[81]));
  AL_DFF_0 al_527fdc5d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[82]));
  AL_DFF_0 al_78b52f9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[83]));
  AL_DFF_0 al_83b9f1b0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[84]));
  AL_DFF_0 al_62ae0238 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[85]));
  AL_DFF_0 al_fd4e3e32 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[86]));
  AL_DFF_0 al_55223ef1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[87]));
  AL_DFF_0 al_f58d59e9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[88]));
  AL_DFF_0 al_97f1c798 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[89]));
  AL_DFF_0 al_5a756331 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[90]));
  AL_DFF_0 al_66037863 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[91]));
  AL_DFF_0 al_d744792c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[92]));
  AL_DFF_0 al_9cd9334b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[93]));
  AL_DFF_0 al_eb160588 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[94]));
  AL_DFF_0 al_e37ea790 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[95]));
  AL_DFF_0 al_a4ffeeed (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[96]));
  AL_DFF_0 al_a83107b6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[97]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[97]));
  AL_DFF_0 al_4a945ba9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[98]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[98]));
  AL_DFF_0 al_b3600540 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[99]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[99]));
  AL_DFF_0 al_ab2d97ea (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[100]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[100]));
  AL_DFF_0 al_210e6643 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[101]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[101]));
  AL_DFF_0 al_90d164d6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[102]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[102]));
  AL_DFF_0 al_a31eebb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[103]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[103]));
  AL_DFF_0 al_f6d95ccf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[104]));
  AL_DFF_0 al_8b87a34 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[105]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[105]));
  AL_DFF_0 al_3f520835 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[106]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[106]));
  AL_DFF_0 al_713c50ec (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[107]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[107]));
  AL_DFF_0 al_a17693b6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[108]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[108]));
  AL_DFF_0 al_a139b7d4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[109]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[109]));
  AL_DFF_0 al_8e2a977a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[110]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[110]));
  AL_DFF_0 al_721a3551 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[111]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[111]));
  AL_DFF_0 al_bb1d80f8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[112]));
  AL_DFF_0 al_10af4d6b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[113]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[113]));
  AL_DFF_0 al_37813ff2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[114]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[114]));
  AL_DFF_0 al_6970c62e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[115]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[115]));
  AL_DFF_0 al_c51045df (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[116]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[116]));
  AL_DFF_0 al_fe42dea0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[117]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[117]));
  AL_DFF_0 al_6ef4165e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[118]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[118]));
  AL_DFF_0 al_6c03c115 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[119]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[119]));
  AL_DFF_0 al_e2555324 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[120]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[120]));
  AL_DFF_0 al_96c50951 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[121]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[121]));
  AL_DFF_0 al_136a99ec (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[122]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[122]));
  AL_DFF_0 al_45273152 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[123]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[123]));
  AL_DFF_0 al_f19222ed (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[124]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[124]));
  AL_DFF_0 al_70ff1c0b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[125]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[125]));
  AL_DFF_0 al_8b5dc73b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[126]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[126]));
  AL_DFF_0 al_edce4d54 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_880499db[127]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32e78cf2[127]));
  AL_DFF_0 al_4b816d6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[0]));
  AL_DFF_0 al_b1d72e39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[3]));
  AL_DFF_0 al_d585493d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[4]));
  AL_DFF_0 al_178ffee3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[5]));
  AL_DFF_0 al_e315b56c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[6]));
  AL_DFF_0 al_cfc32689 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[7]));
  AL_DFF_0 al_aef77eb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[8]));
  AL_DFF_0 al_b2f7ccf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[9]));
  AL_DFF_0 al_78df1793 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[14]));
  AL_DFF_0 al_5592d150 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[15]));
  AL_DFF_0 al_71977513 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[16]));
  AL_DFF_0 al_301d432a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[17]));
  AL_DFF_0 al_6fcc6f41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[18]));
  AL_DFF_0 al_c1fc7b1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[19]));
  AL_DFF_0 al_d9d8811a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[20]));
  AL_DFF_0 al_cd2c9c6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[21]));
  AL_DFF_0 al_8027bfb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[22]));
  AL_DFF_0 al_a5834304 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[23]));
  AL_DFF_0 al_1207b1c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[24]));
  AL_DFF_0 al_cf4bfbc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[25]));
  AL_DFF_0 al_3d08d909 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[26]));
  AL_DFF_0 al_cabe7975 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[27]));
  AL_DFF_0 al_37d0c404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4152494a[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f09d84cf[42]));
  AL_DFF_0 al_986056ef (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[8]));
  AL_DFF_0 al_8e1cee9a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[9]));
  AL_DFF_0 al_1f189370 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[10]));
  AL_DFF_0 al_8fb6cf22 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[11]));
  AL_DFF_0 al_7827dc6d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[12]));
  AL_DFF_0 al_9a383260 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[13]));
  AL_DFF_0 al_bee77bf0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[14]));
  AL_DFF_0 al_cc7ef594 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[15]));
  AL_DFF_0 al_cf94ea74 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[40]));
  AL_DFF_0 al_286de3fb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[41]));
  AL_DFF_0 al_8baf094b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[42]));
  AL_DFF_0 al_8ada06bd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[43]));
  AL_DFF_0 al_5fe6f7d6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[44]));
  AL_DFF_0 al_166cb8ba (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[45]));
  AL_DFF_0 al_594274b5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[46]));
  AL_DFF_0 al_b8bf8c1b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[47]));
  AL_DFF_0 al_44b7ec9a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[72]));
  AL_DFF_0 al_acc59d87 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[73]));
  AL_DFF_0 al_7a78b7bd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[74]));
  AL_DFF_0 al_9a93ae49 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[75]));
  AL_DFF_0 al_6586b59b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[76]));
  AL_DFF_0 al_cad220f4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[77]));
  AL_DFF_0 al_614c6003 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[78]));
  AL_DFF_0 al_171b0d7d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[79]));
  AL_DFF_0 al_73d6e6bc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[104]));
  AL_DFF_0 al_9b1d0ce1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[105]));
  AL_DFF_0 al_e8e5dd74 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[106]));
  AL_DFF_0 al_bbbb4692 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[107]));
  AL_DFF_0 al_6b2f75d2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[108]));
  AL_DFF_0 al_a0e5e08d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[109]));
  AL_DFF_0 al_445828b7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[110]));
  AL_DFF_0 al_6ba45039 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70931fdb[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[111]));
  AL_DFF_0 al_542c83bb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[136]));
  AL_DFF_0 al_5917d439 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[137]));
  AL_DFF_0 al_7f81ed43 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[138]));
  AL_DFF_0 al_b055f1e4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[139]));
  AL_DFF_0 al_bd770059 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[140]));
  AL_DFF_0 al_127a27c0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[141]));
  AL_DFF_0 al_fbd67593 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[142]));
  AL_DFF_0 al_1157f8c9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[143]));
  AL_DFF_0 al_6cef854 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[168]));
  AL_DFF_0 al_f0a8bd1a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[169]));
  AL_DFF_0 al_ad25f68f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[170]));
  AL_DFF_0 al_2d3c48c4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[171]));
  AL_DFF_0 al_c291d5f3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[172]));
  AL_DFF_0 al_38f0239f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[173]));
  AL_DFF_0 al_a394f960 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[174]));
  AL_DFF_0 al_f7ebea43 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[175]));
  AL_DFF_0 al_2500d691 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[200]));
  AL_DFF_0 al_d0c1f672 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[201]));
  AL_DFF_0 al_7c007afe (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[202]));
  AL_DFF_0 al_8d6651a8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[203]));
  AL_DFF_0 al_320a7e03 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[204]));
  AL_DFF_0 al_f4f6a23d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[205]));
  AL_DFF_0 al_7a2c6c9b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[206]));
  AL_DFF_0 al_452f684f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[207]));
  AL_DFF_0 al_5c14a422 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[232]));
  AL_DFF_0 al_5e2c3f1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[233]));
  AL_DFF_0 al_e8129a1f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[234]));
  AL_DFF_0 al_1e0c9cc4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[235]));
  AL_DFF_0 al_d1fb3ba7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[236]));
  AL_DFF_0 al_dcc90faa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[237]));
  AL_DFF_0 al_36318699 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[238]));
  AL_DFF_0 al_95c0f947 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[239]));
  AL_DFF_0 al_64dde9b3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[64]));
  AL_DFF_0 al_8f67f315 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[65]));
  AL_DFF_0 al_50edda47 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[66]));
  AL_DFF_0 al_d2d2bdaf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[67]));
  AL_DFF_0 al_ea9a00aa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[68]));
  AL_DFF_0 al_4184c9b9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[69]));
  AL_DFF_0 al_9f70882c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[70]));
  AL_DFF_0 al_3f5379bd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[71]));
  AL_DFF_0 al_235b72d4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[72]));
  AL_DFF_0 al_5f9c89bb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[73]));
  AL_DFF_0 al_e9946ef3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[74]));
  AL_DFF_0 al_e661c8a1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[75]));
  AL_DFF_0 al_67888b64 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[76]));
  AL_DFF_0 al_f16e0d41 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[77]));
  AL_DFF_0 al_71b67378 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[78]));
  AL_DFF_0 al_47baba08 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[79]));
  AL_DFF_0 al_1d2edfd3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[80]));
  AL_DFF_0 al_da0e4e57 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[81]));
  AL_DFF_0 al_15545f33 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[82]));
  AL_DFF_0 al_de74c375 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[83]));
  AL_DFF_0 al_751ed315 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[84]));
  AL_DFF_0 al_7e9994e7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[85]));
  AL_DFF_0 al_818fb150 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[86]));
  AL_DFF_0 al_7729d7fe (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[87]));
  AL_DFF_0 al_6faa77e1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[88]));
  AL_DFF_0 al_410b4a99 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[89]));
  AL_DFF_0 al_bc5e31ef (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[90]));
  AL_DFF_0 al_3590dfe1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[91]));
  AL_DFF_0 al_e28f2f23 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[92]));
  AL_DFF_0 al_3cc7456a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[93]));
  AL_DFF_0 al_6463792c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[94]));
  AL_DFF_0 al_40ac44ae (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[95]));
  AL_DFF_0 al_4cae7bee (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[96]));
  AL_DFF_0 al_7e237f58 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[97]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[97]));
  AL_DFF_0 al_f06815db (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[98]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[98]));
  AL_DFF_0 al_4146cf96 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[99]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[99]));
  AL_DFF_0 al_aa979f5a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[100]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[100]));
  AL_DFF_0 al_e70a4f39 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[101]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[101]));
  AL_DFF_0 al_c594b6b5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[102]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[102]));
  AL_DFF_0 al_3758ae9a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[103]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[103]));
  AL_DFF_0 al_f648e368 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[104]));
  AL_DFF_0 al_11571e26 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[105]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[105]));
  AL_DFF_0 al_ed7d1dab (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[106]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[106]));
  AL_DFF_0 al_39de41c0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[107]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[107]));
  AL_DFF_0 al_3b0cbe18 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[108]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[108]));
  AL_DFF_0 al_fb5ea3ab (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[109]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[109]));
  AL_DFF_0 al_5113725d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[110]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[110]));
  AL_DFF_0 al_89345b29 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[111]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[111]));
  AL_DFF_0 al_997fef2f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[112]));
  AL_DFF_0 al_1a330b9a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[113]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[113]));
  AL_DFF_0 al_afd11f21 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[114]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[114]));
  AL_DFF_0 al_e3d016a3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[115]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[115]));
  AL_DFF_0 al_17f01b25 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[116]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[116]));
  AL_DFF_0 al_ee786a12 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[117]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[117]));
  AL_DFF_0 al_3921c096 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[118]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[118]));
  AL_DFF_0 al_e535ba41 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[119]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[119]));
  AL_DFF_0 al_10bfc528 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[120]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[120]));
  AL_DFF_0 al_6a5141a8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[121]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[121]));
  AL_DFF_0 al_b7a354b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[122]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[122]));
  AL_DFF_0 al_76827e7b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[123]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[123]));
  AL_DFF_0 al_7ffeee00 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[124]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[124]));
  AL_DFF_0 al_613ebdfa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[125]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[125]));
  AL_DFF_0 al_a23bda7d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[126]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[126]));
  AL_DFF_0 al_a6c2610f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2982a0b8[127]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70931fdb[127]));
  AL_DFF_0 al_1097f80d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[16]));
  AL_DFF_0 al_94c7308c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[17]));
  AL_DFF_0 al_4ceb8d33 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[18]));
  AL_DFF_0 al_4a42af80 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[19]));
  AL_DFF_0 al_d65c8eb5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[20]));
  AL_DFF_0 al_e8653f92 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[21]));
  AL_DFF_0 al_9a357cdf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[22]));
  AL_DFF_0 al_13ea8e96 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[23]));
  AL_DFF_0 al_6876a074 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[48]));
  AL_DFF_0 al_b03fce5c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[49]));
  AL_DFF_0 al_c4969076 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[50]));
  AL_DFF_0 al_d673b585 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[51]));
  AL_DFF_0 al_1a9f553f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[52]));
  AL_DFF_0 al_9b9a143b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[53]));
  AL_DFF_0 al_e27d7c1a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[54]));
  AL_DFF_0 al_5ddb7350 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[55]));
  AL_DFF_0 al_220e1a60 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[80]));
  AL_DFF_0 al_a5c42120 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[81]));
  AL_DFF_0 al_4d70f27e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[82]));
  AL_DFF_0 al_e77e7a9f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[83]));
  AL_DFF_0 al_4357ea26 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[84]));
  AL_DFF_0 al_bcf2e69d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[85]));
  AL_DFF_0 al_d7a8b2c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[86]));
  AL_DFF_0 al_29d9f13e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[87]));
  AL_DFF_0 al_2fea0b1f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[112]));
  AL_DFF_0 al_385d83ac (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[113]));
  AL_DFF_0 al_2815fedf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[114]));
  AL_DFF_0 al_e24f4c57 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[115]));
  AL_DFF_0 al_4675e78c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[116]));
  AL_DFF_0 al_87ab5114 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[117]));
  AL_DFF_0 al_51e1996e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[118]));
  AL_DFF_0 al_6c2f0b95 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3f231cd[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[119]));
  AL_DFF_0 al_764d4698 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[144]));
  AL_DFF_0 al_f612b691 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[145]));
  AL_DFF_0 al_ff24389a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[146]));
  AL_DFF_0 al_5b944e54 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[147]));
  AL_DFF_0 al_13c39bcf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[148]));
  AL_DFF_0 al_8dd43e10 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[149]));
  AL_DFF_0 al_f41e61dd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[150]));
  AL_DFF_0 al_df01ad70 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[151]));
  AL_DFF_0 al_2ee2d688 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[176]));
  AL_DFF_0 al_e1212c85 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[177]));
  AL_DFF_0 al_39fd445b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[178]));
  AL_DFF_0 al_ff392724 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[179]));
  AL_DFF_0 al_d835c3f8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[180]));
  AL_DFF_0 al_854a7c7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[181]));
  AL_DFF_0 al_bd9d023f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[182]));
  AL_DFF_0 al_b16cc0dd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[183]));
  AL_DFF_0 al_c4ca6f80 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[208]));
  AL_DFF_0 al_e74d712a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[209]));
  AL_DFF_0 al_14b3fcd2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[210]));
  AL_DFF_0 al_8fac4846 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[211]));
  AL_DFF_0 al_21a67a7e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[212]));
  AL_DFF_0 al_74129af4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[213]));
  AL_DFF_0 al_b7bec9a8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[214]));
  AL_DFF_0 al_aa610e4b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[215]));
  AL_DFF_0 al_18f190dc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[240]));
  AL_DFF_0 al_238e10e2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[241]));
  AL_DFF_0 al_bba45236 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[242]));
  AL_DFF_0 al_699efb5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[243]));
  AL_DFF_0 al_61f943be (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[244]));
  AL_DFF_0 al_bad300e5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[245]));
  AL_DFF_0 al_24f968b8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[246]));
  AL_DFF_0 al_eb51dab8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[247]));
  AL_DFF_0 al_e08fc2e6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[64]));
  AL_DFF_0 al_b801517c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[65]));
  AL_DFF_0 al_ad6e0739 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[66]));
  AL_DFF_0 al_ee76b37d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[67]));
  AL_DFF_0 al_342eb35e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[68]));
  AL_DFF_0 al_485ae57b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[69]));
  AL_DFF_0 al_4dfb97c6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[70]));
  AL_DFF_0 al_d3c917e3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[71]));
  AL_DFF_0 al_aa48f78 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[72]));
  AL_DFF_0 al_3b0f05eb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[73]));
  AL_DFF_0 al_e6f32036 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[74]));
  AL_DFF_0 al_fe2dd327 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[75]));
  AL_DFF_0 al_cc537149 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[76]));
  AL_DFF_0 al_276b6cb4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[77]));
  AL_DFF_0 al_ebfb1bab (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[78]));
  AL_DFF_0 al_aa6a7c5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[79]));
  AL_DFF_0 al_f15c0cf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[80]));
  AL_DFF_0 al_3196cd3f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[81]));
  AL_DFF_0 al_51d8da7b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[82]));
  AL_DFF_0 al_148f2be (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[83]));
  AL_DFF_0 al_fe20a5d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[84]));
  AL_DFF_0 al_13048c5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[85]));
  AL_DFF_0 al_86159169 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[86]));
  AL_DFF_0 al_a828d9c1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[87]));
  AL_DFF_0 al_4f6ea3d6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[88]));
  AL_DFF_0 al_f592dd6e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[89]));
  AL_DFF_0 al_b64d231d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[90]));
  AL_DFF_0 al_630ab698 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[91]));
  AL_DFF_0 al_bc54a9e2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[92]));
  AL_DFF_0 al_b38c2157 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[93]));
  AL_DFF_0 al_3ddc5af0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[94]));
  AL_DFF_0 al_7ddf7c79 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[95]));
  AL_DFF_0 al_621e4232 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[96]));
  AL_DFF_0 al_c7ff1e53 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[97]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[97]));
  AL_DFF_0 al_79a0cdff (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[98]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[98]));
  AL_DFF_0 al_d327f4e7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[99]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[99]));
  AL_DFF_0 al_afdc5307 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[100]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[100]));
  AL_DFF_0 al_d2bf4da9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[101]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[101]));
  AL_DFF_0 al_3e563f06 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[102]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[102]));
  AL_DFF_0 al_41bbc52e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[103]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[103]));
  AL_DFF_0 al_113c1af7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[104]));
  AL_DFF_0 al_d0835c86 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[105]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[105]));
  AL_DFF_0 al_aa4228c1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[106]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[106]));
  AL_DFF_0 al_c032ec60 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[107]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[107]));
  AL_DFF_0 al_8962fcb3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[108]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[108]));
  AL_DFF_0 al_2c0e4d92 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[109]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[109]));
  AL_DFF_0 al_58cf4fca (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[110]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[110]));
  AL_DFF_0 al_6df3734e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[111]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[111]));
  AL_DFF_0 al_a84df3db (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[112]));
  AL_DFF_0 al_57f12c73 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[113]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[113]));
  AL_DFF_0 al_2634616a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[114]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[114]));
  AL_DFF_0 al_1e3dd70f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[115]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[115]));
  AL_DFF_0 al_4e747336 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[116]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[116]));
  AL_DFF_0 al_32d935a9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[117]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[117]));
  AL_DFF_0 al_487a3aae (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[118]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[118]));
  AL_DFF_0 al_6630d3a7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[119]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[119]));
  AL_DFF_0 al_97398806 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[120]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[120]));
  AL_DFF_0 al_34575485 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[121]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[121]));
  AL_DFF_0 al_7a5c5453 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[122]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[122]));
  AL_DFF_0 al_eb6bb407 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[123]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[123]));
  AL_DFF_0 al_c94e15c5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[124]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[124]));
  AL_DFF_0 al_5238a398 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[125]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[125]));
  AL_DFF_0 al_2321936e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[126]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[126]));
  AL_DFF_0 al_4456c2d5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cde313f8[127]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3f231cd[127]));
  AL_DFF_0 al_81c53c21 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[24]));
  AL_DFF_0 al_dc10de62 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[25]));
  AL_DFF_0 al_4422bb01 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[26]));
  AL_DFF_0 al_2f918bda (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[27]));
  AL_DFF_0 al_6af95287 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[28]));
  AL_DFF_0 al_536bf424 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[29]));
  AL_DFF_0 al_62ae4625 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[30]));
  AL_DFF_0 al_221a223e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[31]));
  AL_DFF_0 al_81d47a49 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[56]));
  AL_DFF_0 al_d36418e4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[57]));
  AL_DFF_0 al_b5342725 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[58]));
  AL_DFF_0 al_be149785 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[59]));
  AL_DFF_0 al_6e7b37cf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[60]));
  AL_DFF_0 al_41bd806c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[61]));
  AL_DFF_0 al_9c03134d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[62]));
  AL_DFF_0 al_2072993 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[63]));
  AL_DFF_0 al_4063a623 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[88]));
  AL_DFF_0 al_dd9874cf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[89]));
  AL_DFF_0 al_3825a735 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[90]));
  AL_DFF_0 al_95f5aae9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[91]));
  AL_DFF_0 al_2f0f63aa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[92]));
  AL_DFF_0 al_8893030a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[93]));
  AL_DFF_0 al_f44fd44c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[94]));
  AL_DFF_0 al_3a15483b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[95]));
  AL_DFF_0 al_aefe6e97 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[120]));
  AL_DFF_0 al_b3918134 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[121]));
  AL_DFF_0 al_ca2ef8f3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[122]));
  AL_DFF_0 al_462d6e97 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[123]));
  AL_DFF_0 al_c83d1757 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[124]));
  AL_DFF_0 al_270d7dd2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[125]));
  AL_DFF_0 al_683d5bf8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[126]));
  AL_DFF_0 al_77a0b877 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1c5f121[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[127]));
  AL_DFF_0 al_319d5d3c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[152]));
  AL_DFF_0 al_fcfffd73 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[153]));
  AL_DFF_0 al_f5063791 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[154]));
  AL_DFF_0 al_7de751bb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[155]));
  AL_DFF_0 al_320858b1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[156]));
  AL_DFF_0 al_25534dfe (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[157]));
  AL_DFF_0 al_db4a93eb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[158]));
  AL_DFF_0 al_f045cdd1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[159]));
  AL_DFF_0 al_a8564742 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[184]));
  AL_DFF_0 al_9bb588e3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[185]));
  AL_DFF_0 al_3865cd88 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[186]));
  AL_DFF_0 al_8b8e9da8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[187]));
  AL_DFF_0 al_e4d6497e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[188]));
  AL_DFF_0 al_a7e672b3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[189]));
  AL_DFF_0 al_10ca311 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[190]));
  AL_DFF_0 al_3234ef58 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[191]));
  AL_DFF_0 al_84d47648 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[216]));
  AL_DFF_0 al_dff26d57 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[217]));
  AL_DFF_0 al_3e9cb2bd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[218]));
  AL_DFF_0 al_6946a36 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[219]));
  AL_DFF_0 al_dfb4355e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[220]));
  AL_DFF_0 al_903d0989 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[221]));
  AL_DFF_0 al_28749056 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[222]));
  AL_DFF_0 al_321fda2c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[223]));
  AL_DFF_0 al_1515197d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[248]));
  AL_DFF_0 al_a6ad272e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[249]));
  AL_DFF_0 al_71e8faf2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[250]));
  AL_DFF_0 al_b1a3ebc1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[251]));
  AL_DFF_0 al_e0b59554 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[252]));
  AL_DFF_0 al_729276d8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[253]));
  AL_DFF_0 al_bb558dec (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[254]));
  AL_DFF_0 al_7ad52952 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_p[255]));
  AL_DFF_0 al_4b563662 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[64]));
  AL_DFF_0 al_99518d37 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[65]));
  AL_DFF_0 al_444149bb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[66]));
  AL_DFF_0 al_c35a7709 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[67]));
  AL_DFF_0 al_1d77b154 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[68]));
  AL_DFF_0 al_e529c437 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[69]));
  AL_DFF_0 al_c472253b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[70]));
  AL_DFF_0 al_e0cd2b9f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[71]));
  AL_DFF_0 al_b6c3bfcd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[72]));
  AL_DFF_0 al_de5bd38d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[73]));
  AL_DFF_0 al_8215b03 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[74]));
  AL_DFF_0 al_e0ce2612 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[75]));
  AL_DFF_0 al_22586825 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[76]));
  AL_DFF_0 al_f80fbc48 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[77]));
  AL_DFF_0 al_2600e527 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[78]));
  AL_DFF_0 al_9af7a21d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[79]));
  AL_DFF_0 al_fcdb658e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[80]));
  AL_DFF_0 al_9c873833 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[81]));
  AL_DFF_0 al_5c987dd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[82]));
  AL_DFF_0 al_ad047ded (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[83]));
  AL_DFF_0 al_c6ae0da9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[84]));
  AL_DFF_0 al_75474ae3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[85]));
  AL_DFF_0 al_6e68e8d9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[86]));
  AL_DFF_0 al_876a5fb6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[87]));
  AL_DFF_0 al_e366920b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[88]));
  AL_DFF_0 al_f9f6a35f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[89]));
  AL_DFF_0 al_44b2ad80 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[90]));
  AL_DFF_0 al_7fa4f7da (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[91]));
  AL_DFF_0 al_b4f3d9ae (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[92]));
  AL_DFF_0 al_821f42d3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[93]));
  AL_DFF_0 al_65211d1a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[94]));
  AL_DFF_0 al_b336834a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[95]));
  AL_DFF_0 al_e11ffefc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[96]));
  AL_DFF_0 al_177a1a5d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[97]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[97]));
  AL_DFF_0 al_4fb68726 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[98]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[98]));
  AL_DFF_0 al_6f82bc0c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[99]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[99]));
  AL_DFF_0 al_26b8563c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[100]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[100]));
  AL_DFF_0 al_54fc95ee (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[101]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[101]));
  AL_DFF_0 al_49763460 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[102]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[102]));
  AL_DFF_0 al_6bac58c0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[103]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[103]));
  AL_DFF_0 al_9ec22f41 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[104]));
  AL_DFF_0 al_f14e7ec4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[105]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[105]));
  AL_DFF_0 al_8bb66261 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[106]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[106]));
  AL_DFF_0 al_84c22b28 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[107]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[107]));
  AL_DFF_0 al_82834e5e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[108]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[108]));
  AL_DFF_0 al_557ac978 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[109]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[109]));
  AL_DFF_0 al_b4988127 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[110]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[110]));
  AL_DFF_0 al_b7cefd4a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[111]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[111]));
  AL_DFF_0 al_a2c3c3e8 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[112]));
  AL_DFF_0 al_e2ae887f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[113]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[113]));
  AL_DFF_0 al_f5d5535e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[114]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[114]));
  AL_DFF_0 al_fc6d05b7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[115]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[115]));
  AL_DFF_0 al_235c93a9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[116]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[116]));
  AL_DFF_0 al_bed02244 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[117]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[117]));
  AL_DFF_0 al_fc4fdd7f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[118]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[118]));
  AL_DFF_0 al_43879ee1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[119]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[119]));
  AL_DFF_0 al_22467619 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[120]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[120]));
  AL_DFF_0 al_aa8104e9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[121]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[121]));
  AL_DFF_0 al_a5cffed1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[122]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[122]));
  AL_DFF_0 al_bf352905 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[123]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[123]));
  AL_DFF_0 al_75a71721 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[124]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[124]));
  AL_DFF_0 al_762abea0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[125]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[125]));
  AL_DFF_0 al_ff3a5fe6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[126]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[126]));
  AL_DFF_0 al_37d6fafd (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b43737f6[127]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1c5f121[127]));
  AL_DFF_0 al_bfab052e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef9accde),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cc4d831c[0]));
  AL_DFF_0 al_9777964c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cc4d831c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cc4d831c[1]));
  AL_DFF_0 al_35718646 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cc4d831c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f7c5f81));
  AL_DFF_0 al_3b57c4b1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8679dfa[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8679dfa[0]));
  AL_DFF_0 al_c423050c (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8679dfa[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8679dfa[3]));
  AL_DFF_0 al_8aa9333a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea19deeb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8679dfa[4]));
  AL_DFF_0 al_b60926ae (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80aa352a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8679dfa[7]));
  AL_DFF_0 al_e2adfe2a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea19deeb[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8679dfa[8]));
  AL_DFF_0 al_e0896cab (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4340e4e7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[0]));
  AL_DFF_0 al_b634f8aa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4340e4e7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[4]));
  AL_DFF_0 al_641771bc (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4340e4e7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[8]));
  AL_DFF_0 al_f39a0619 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4340e4e7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[12]));
  AL_DFF_0 al_c01eaf5f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[16]));
  AL_DFF_0 al_2e44442a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[20]));
  AL_DFF_0 al_1c0658e5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[24]));
  AL_DFF_0 al_248889fb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[28]));
  AL_DFF_0 al_d6a35e4f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4340e4e7[8]));
  AL_DFF_0 al_9c88b4e2 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4340e4e7[9]));
  AL_DFF_0 al_464b3345 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4340e4e7[10]));
  AL_DFF_0 al_165ac4ed (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4340e4e7[11]));
  AL_DFF_0 al_2a76fc66 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4340e4e7[12]));
  AL_DFF_0 al_d26b7a13 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4340e4e7[13]));
  AL_DFF_0 al_bf378c39 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4340e4e7[14]));
  AL_DFF_0 al_9e889178 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_523e9f7a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4340e4e7[15]));
  AL_DFF_0 al_da563af6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55ed1bfd[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[1]));
  AL_DFF_0 al_6456f60e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55ed1bfd[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[5]));
  AL_DFF_0 al_1fc3d067 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55ed1bfd[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[9]));
  AL_DFF_0 al_d183d9e1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55ed1bfd[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[13]));
  AL_DFF_0 al_abfb23f6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[17]));
  AL_DFF_0 al_a5715c21 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[21]));
  AL_DFF_0 al_7c432a0d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[25]));
  AL_DFF_0 al_c6d2c12f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[29]));
  AL_DFF_0 al_bf4568e1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ed1bfd[8]));
  AL_DFF_0 al_1cbadba7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ed1bfd[9]));
  AL_DFF_0 al_7efcef09 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ed1bfd[10]));
  AL_DFF_0 al_885b0dbf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ed1bfd[11]));
  AL_DFF_0 al_eece5b47 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ed1bfd[12]));
  AL_DFF_0 al_6395d0d7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ed1bfd[13]));
  AL_DFF_0 al_d719992f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ed1bfd[14]));
  AL_DFF_0 al_18cc4360 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ef9bc8c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ed1bfd[15]));
  AL_DFF_0 al_2999d99d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0d99cb1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[2]));
  AL_DFF_0 al_ceaafa9b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0d99cb1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[6]));
  AL_DFF_0 al_5b342b9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0d99cb1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[10]));
  AL_DFF_0 al_af6c52e0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0d99cb1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[14]));
  AL_DFF_0 al_611e7590 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[18]));
  AL_DFF_0 al_4b947abf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[22]));
  AL_DFF_0 al_d886403a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[26]));
  AL_DFF_0 al_b0db8c6b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[30]));
  AL_DFF_0 al_41169092 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0d99cb1[8]));
  AL_DFF_0 al_790642f0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0d99cb1[9]));
  AL_DFF_0 al_104cb45f (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0d99cb1[10]));
  AL_DFF_0 al_fa90ad2e (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0d99cb1[11]));
  AL_DFF_0 al_a7877fdb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0d99cb1[12]));
  AL_DFF_0 al_befb7426 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0d99cb1[13]));
  AL_DFF_0 al_2248c631 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0d99cb1[14]));
  AL_DFF_0 al_da6963a6 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1aabbd4[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0d99cb1[15]));
  AL_DFF_0 al_d3240989 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f949a7ee[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[3]));
  AL_DFF_0 al_b910f1b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f949a7ee[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[7]));
  AL_DFF_0 al_52f043fa (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f949a7ee[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[11]));
  AL_DFF_0 al_d2eaf820 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f949a7ee[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[15]));
  AL_DFF_0 al_35f1797b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[19]));
  AL_DFF_0 al_1c9522f0 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[23]));
  AL_DFF_0 al_51448ff9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[27]));
  AL_DFF_0 al_2c134ad4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_wrdata_mask_p[31]));
  AL_DFF_0 al_1bc1b851 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f949a7ee[8]));
  AL_DFF_0 al_e84591e1 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f949a7ee[9]));
  AL_DFF_0 al_38f8b2fb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f949a7ee[10]));
  AL_DFF_0 al_c0e93a01 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f949a7ee[11]));
  AL_DFF_0 al_38f5da28 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f949a7ee[12]));
  AL_DFF_0 al_f3774a53 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f949a7ee[13]));
  AL_DFF_0 al_955db465 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f949a7ee[14]));
  AL_DFF_0 al_81358d8a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f2a09ff[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f949a7ee[15]));
  AL_DFF_0 al_5bcb5922 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_95504971[136]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[0]));
  AL_DFF_0 al_8e3c4e97 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_95504971[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[3]));
  AL_DFF_0 al_6290b23a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_95504971[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[4]));
  AL_DFF_0 al_2852a1f7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_95504971[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[5]));
  AL_DFF_0 al_d7abc4de (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_95504971[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[6]));
  AL_DFF_0 al_50c4444b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_95504971[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[7]));
  AL_DFF_0 al_799aacce (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_95504971[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[8]));
  AL_DFF_0 al_91fc80d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_95504971[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[9]));
  AL_DFF_0 al_eeb58902 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eb9aa630[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[14]));
  AL_DFF_0 al_248d87b9 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_534b111d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[15]));
  AL_DFF_0 al_9da9738a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_39691102[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[16]));
  AL_DFF_0 al_f35225b5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_304bc4cf[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[17]));
  AL_DFF_0 al_12c71870 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_421a630e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[18]));
  AL_DFF_0 al_fb4d1caf (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2cee9b7b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[19]));
  AL_DFF_0 al_421fd850 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2f77b9ea[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[20]));
  AL_DFF_0 al_f35ab210 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7a66cc8[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[21]));
  AL_DFF_0 al_9070903d (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bce3182d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[22]));
  AL_DFF_0 al_d60adf00 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_636a0d93[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[23]));
  AL_DFF_0 al_7702dae (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3c0a4ef0[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[24]));
  AL_DFF_0 al_ff1841b5 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ecc8e317[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[25]));
  AL_DFF_0 al_73fa064b (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c8b553c9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[26]));
  AL_DFF_0 al_2316afdb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_92812db2[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[27]));
  AL_DFF_0 al_cb96c328 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eb9aa630[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4152494a[42]));
  AL_DFF_0 al_c5dce424 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[0]));
  AL_DFF_0 al_864b4542 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[1]));
  AL_DFF_0 al_5155dc64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[2]));
  AL_DFF_0 al_c320b404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[3]));
  AL_DFF_0 al_9a4813ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[4]));
  AL_DFF_0 al_86a5cc3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[5]));
  AL_DFF_0 al_ed71e768 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[9]));
  AL_DFF_0 al_73a03bc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[10]));
  AL_DFF_0 al_b5584a0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80bec816[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dfi_bank_p[11]));
  AL_DFF_0 al_3962c670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[0]));
  AL_DFF_0 al_a0731c19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[1]));
  AL_DFF_0 al_eccf7dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[2]));
  AL_DFF_0 al_e4069183 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[3]));
  AL_DFF_0 al_4d817956 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[4]));
  AL_DFF_0 al_5bf6abf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[5]));
  AL_DFF_0 al_c9504670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[9]));
  AL_DFF_0 al_4db74a54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[10]));
  AL_DFF_0 al_348cdb3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b678b52[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80bec816[11]));
  AL_DFF_0 al_bfdc6ba (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3639d7e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[0]));
  AL_DFF_0 al_453fefc7 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_18fbbb0f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[1]));
  AL_DFF_0 al_737c7128 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_779bd70c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[2]));
  AL_DFF_0 al_4175a3a3 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3639d7e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[3]));
  AL_DFF_0 al_e06b0df4 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_18fbbb0f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[4]));
  AL_DFF_0 al_45417c1a (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_779bd70c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[5]));
  AL_DFF_0 al_2355cdbb (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3639d7e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[9]));
  AL_DFF_0 al_bd9cef13 (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_18fbbb0f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[10]));
  AL_DFF_0 al_5bfe0df (
    .ar(rst),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_779bd70c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b678b52[11]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_ae6c656 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[84]),
    .e(al_3e0d53ab[100]),
    .o(al_2982a0b8[100]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c25d4c39 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[85]),
    .e(al_3e0d53ab[101]),
    .o(al_2982a0b8[101]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_8c4f7fc6 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[86]),
    .e(al_3e0d53ab[102]),
    .o(al_2982a0b8[102]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_303271cd (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[87]),
    .e(al_3e0d53ab[103]),
    .o(al_2982a0b8[103]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_f78496d5 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[88]),
    .e(al_3e0d53ab[104]),
    .o(al_2982a0b8[104]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_8b4d1bec (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[89]),
    .e(al_3e0d53ab[105]),
    .o(al_2982a0b8[105]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_da76e40f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[90]),
    .e(al_3e0d53ab[106]),
    .o(al_2982a0b8[106]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_8b4ad0a6 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[91]),
    .e(al_3e0d53ab[107]),
    .o(al_2982a0b8[107]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_569c1dfd (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[92]),
    .e(al_3e0d53ab[108]),
    .o(al_2982a0b8[108]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_1133bbe7 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[93]),
    .e(al_3e0d53ab[109]),
    .o(al_2982a0b8[109]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_560cee68 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[94]),
    .e(al_3e0d53ab[110]),
    .o(al_2982a0b8[110]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_d4846b29 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[95]),
    .e(al_3e0d53ab[111]),
    .o(al_2982a0b8[111]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_4f7ac13f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[96]),
    .e(al_3e0d53ab[112]),
    .o(al_2982a0b8[112]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_316322a7 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[97]),
    .e(al_3e0d53ab[113]),
    .o(al_2982a0b8[113]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c0cbe362 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[98]),
    .e(al_3e0d53ab[114]),
    .o(al_2982a0b8[114]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_be0d4e3 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[99]),
    .e(al_3e0d53ab[115]),
    .o(al_2982a0b8[115]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_8d03f4be (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[100]),
    .e(al_3e0d53ab[116]),
    .o(al_2982a0b8[116]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_8631f1a7 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[101]),
    .e(al_3e0d53ab[117]),
    .o(al_2982a0b8[117]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_5330d79f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[102]),
    .e(al_3e0d53ab[118]),
    .o(al_2982a0b8[118]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c1443acf (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[103]),
    .e(al_3e0d53ab[119]),
    .o(al_2982a0b8[119]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_4593f56f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[104]),
    .e(al_3e0d53ab[120]),
    .o(al_2982a0b8[120]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_f9939639 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[105]),
    .e(al_3e0d53ab[121]),
    .o(al_2982a0b8[121]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_203fea0d (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[106]),
    .e(al_3e0d53ab[122]),
    .o(al_2982a0b8[122]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_9795498e (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[107]),
    .e(al_3e0d53ab[123]),
    .o(al_2982a0b8[123]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_aa87e996 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[108]),
    .e(al_3e0d53ab[124]),
    .o(al_2982a0b8[124]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_94e317d9 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[109]),
    .e(al_3e0d53ab[125]),
    .o(al_2982a0b8[125]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_bc3e128d (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[110]),
    .e(al_3e0d53ab[126]),
    .o(al_2982a0b8[126]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_f20866c (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[111]),
    .e(al_3e0d53ab[127]),
    .o(al_2982a0b8[127]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_e1a71db2 (
    .a(al_25e28b94),
    .b(al_70931fdb[96]),
    .c(al_3e0d53ab[64]),
    .o(al_2982a0b8[32]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_6b6fe5bd (
    .a(al_25e28b94),
    .b(al_70931fdb[97]),
    .c(al_3e0d53ab[65]),
    .o(al_2982a0b8[33]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_afb8b4fd (
    .a(al_25e28b94),
    .b(al_70931fdb[98]),
    .c(al_3e0d53ab[66]),
    .o(al_2982a0b8[34]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_b1360d26 (
    .a(al_25e28b94),
    .b(al_70931fdb[99]),
    .c(al_3e0d53ab[67]),
    .o(al_2982a0b8[35]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_dd747053 (
    .a(al_25e28b94),
    .b(al_70931fdb[100]),
    .c(al_3e0d53ab[68]),
    .o(al_2982a0b8[36]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_4790cbad (
    .a(al_25e28b94),
    .b(al_70931fdb[101]),
    .c(al_3e0d53ab[69]),
    .o(al_2982a0b8[37]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_c601c3f3 (
    .a(al_25e28b94),
    .b(al_70931fdb[102]),
    .c(al_3e0d53ab[70]),
    .o(al_2982a0b8[38]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9869a76f (
    .a(al_25e28b94),
    .b(al_70931fdb[103]),
    .c(al_3e0d53ab[71]),
    .o(al_2982a0b8[39]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_ff152b17 (
    .a(al_25e28b94),
    .b(al_70931fdb[104]),
    .c(al_3e0d53ab[72]),
    .o(al_2982a0b8[40]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_5a402d9f (
    .a(al_25e28b94),
    .b(al_70931fdb[105]),
    .c(al_3e0d53ab[73]),
    .o(al_2982a0b8[41]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9e92239d (
    .a(al_25e28b94),
    .b(al_70931fdb[106]),
    .c(al_3e0d53ab[74]),
    .o(al_2982a0b8[42]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9a2e3364 (
    .a(al_25e28b94),
    .b(al_70931fdb[107]),
    .c(al_3e0d53ab[75]),
    .o(al_2982a0b8[43]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_5bcabe6d (
    .a(al_25e28b94),
    .b(al_70931fdb[108]),
    .c(al_3e0d53ab[76]),
    .o(al_2982a0b8[44]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_87d3571d (
    .a(al_25e28b94),
    .b(al_70931fdb[109]),
    .c(al_3e0d53ab[77]),
    .o(al_2982a0b8[45]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_5e7c2001 (
    .a(al_25e28b94),
    .b(al_70931fdb[110]),
    .c(al_3e0d53ab[78]),
    .o(al_2982a0b8[46]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_d885f0b1 (
    .a(al_25e28b94),
    .b(al_70931fdb[111]),
    .c(al_3e0d53ab[79]),
    .o(al_2982a0b8[47]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_bfdd5198 (
    .a(al_25e28b94),
    .b(al_70931fdb[112]),
    .c(al_3e0d53ab[80]),
    .o(al_2982a0b8[48]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_da2cca98 (
    .a(al_25e28b94),
    .b(al_70931fdb[113]),
    .c(al_3e0d53ab[81]),
    .o(al_2982a0b8[49]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_c29b7790 (
    .a(al_25e28b94),
    .b(al_70931fdb[114]),
    .c(al_3e0d53ab[82]),
    .o(al_2982a0b8[50]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_798cdd13 (
    .a(al_25e28b94),
    .b(al_70931fdb[115]),
    .c(al_3e0d53ab[83]),
    .o(al_2982a0b8[51]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_5b6bd946 (
    .a(al_25e28b94),
    .b(al_70931fdb[116]),
    .c(al_3e0d53ab[84]),
    .o(al_2982a0b8[52]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_f34a3639 (
    .a(al_25e28b94),
    .b(al_70931fdb[117]),
    .c(al_3e0d53ab[85]),
    .o(al_2982a0b8[53]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_4743201e (
    .a(al_25e28b94),
    .b(al_70931fdb[118]),
    .c(al_3e0d53ab[86]),
    .o(al_2982a0b8[54]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_97c993ff (
    .a(al_25e28b94),
    .b(al_70931fdb[119]),
    .c(al_3e0d53ab[87]),
    .o(al_2982a0b8[55]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_1cf30d99 (
    .a(al_25e28b94),
    .b(al_70931fdb[120]),
    .c(al_3e0d53ab[88]),
    .o(al_2982a0b8[56]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_aec2efcc (
    .a(al_25e28b94),
    .b(al_70931fdb[121]),
    .c(al_3e0d53ab[89]),
    .o(al_2982a0b8[57]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_d2db4df2 (
    .a(al_25e28b94),
    .b(al_70931fdb[122]),
    .c(al_3e0d53ab[90]),
    .o(al_2982a0b8[58]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_a5b6bced (
    .a(al_25e28b94),
    .b(al_70931fdb[123]),
    .c(al_3e0d53ab[91]),
    .o(al_2982a0b8[59]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_66e935cc (
    .a(al_25e28b94),
    .b(al_70931fdb[124]),
    .c(al_3e0d53ab[92]),
    .o(al_2982a0b8[60]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_60eaab35 (
    .a(al_25e28b94),
    .b(al_70931fdb[125]),
    .c(al_3e0d53ab[93]),
    .o(al_2982a0b8[61]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_d1e96c90 (
    .a(al_25e28b94),
    .b(al_70931fdb[126]),
    .c(al_3e0d53ab[94]),
    .o(al_2982a0b8[62]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_11890c1c (
    .a(al_25e28b94),
    .b(al_70931fdb[127]),
    .c(al_3e0d53ab[95]),
    .o(al_2982a0b8[63]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_4f6deef7 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[64]),
    .e(al_3e0d53ab[96]),
    .o(al_2982a0b8[64]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_448cae0b (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[65]),
    .e(al_3e0d53ab[97]),
    .o(al_2982a0b8[65]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_876a11e6 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[66]),
    .e(al_3e0d53ab[98]),
    .o(al_2982a0b8[66]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_63fe51e4 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[67]),
    .e(al_3e0d53ab[99]),
    .o(al_2982a0b8[67]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_c386d068 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[68]),
    .e(al_3e0d53ab[100]),
    .o(al_2982a0b8[68]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_c8545477 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[69]),
    .e(al_3e0d53ab[101]),
    .o(al_2982a0b8[69]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_c0101ff2 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[70]),
    .e(al_3e0d53ab[102]),
    .o(al_2982a0b8[70]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_6fcb38ef (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[71]),
    .e(al_3e0d53ab[103]),
    .o(al_2982a0b8[71]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_4e88c896 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[72]),
    .e(al_3e0d53ab[104]),
    .o(al_2982a0b8[72]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_8c669465 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[73]),
    .e(al_3e0d53ab[105]),
    .o(al_2982a0b8[73]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_6cb1ff71 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[74]),
    .e(al_3e0d53ab[106]),
    .o(al_2982a0b8[74]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_b83595cb (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[75]),
    .e(al_3e0d53ab[107]),
    .o(al_2982a0b8[75]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_aaa633cc (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[76]),
    .e(al_3e0d53ab[108]),
    .o(al_2982a0b8[76]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_de6576b8 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[77]),
    .e(al_3e0d53ab[109]),
    .o(al_2982a0b8[77]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_7eb191a9 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[78]),
    .e(al_3e0d53ab[110]),
    .o(al_2982a0b8[78]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_9cb17ac8 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[79]),
    .e(al_3e0d53ab[111]),
    .o(al_2982a0b8[79]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_280ae1d7 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[64]),
    .e(al_3e0d53ab[80]),
    .f(al_3e0d53ab[112]),
    .o(al_84d9df21));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_7590ed12 (
    .a(al_84d9df21),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[80]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_4a3d385a (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[65]),
    .e(al_3e0d53ab[81]),
    .f(al_3e0d53ab[113]),
    .o(al_786e90e));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ccab9345 (
    .a(al_786e90e),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[81]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_d1babdaa (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[66]),
    .e(al_3e0d53ab[82]),
    .f(al_3e0d53ab[114]),
    .o(al_e56639b1));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e75031cf (
    .a(al_e56639b1),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[82]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_9f5a3253 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[67]),
    .e(al_3e0d53ab[83]),
    .f(al_3e0d53ab[115]),
    .o(al_373390f0));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_88022153 (
    .a(al_373390f0),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[83]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_6afb6944 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[68]),
    .e(al_3e0d53ab[84]),
    .f(al_3e0d53ab[116]),
    .o(al_97ed8d08));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6e471f4c (
    .a(al_97ed8d08),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[84]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_acdc7d45 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[69]),
    .e(al_3e0d53ab[85]),
    .f(al_3e0d53ab[117]),
    .o(al_75463750));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_621155ac (
    .a(al_75463750),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[85]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_7ed8e6ee (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[70]),
    .e(al_3e0d53ab[86]),
    .f(al_3e0d53ab[118]),
    .o(al_4124b4b4));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_46742b07 (
    .a(al_4124b4b4),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[86]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_cab30491 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[71]),
    .e(al_3e0d53ab[87]),
    .f(al_3e0d53ab[119]),
    .o(al_202cea3f));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_45829600 (
    .a(al_202cea3f),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[87]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_6ee56929 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[72]),
    .e(al_3e0d53ab[88]),
    .f(al_3e0d53ab[120]),
    .o(al_19d71bde));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_1005fd2 (
    .a(al_19d71bde),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[88]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_4479a6d8 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[73]),
    .e(al_3e0d53ab[89]),
    .f(al_3e0d53ab[121]),
    .o(al_29e00248));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cb3a234d (
    .a(al_29e00248),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[89]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_89e6ba62 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[74]),
    .e(al_3e0d53ab[90]),
    .f(al_3e0d53ab[122]),
    .o(al_f486e5f));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b27cd9e6 (
    .a(al_f486e5f),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[90]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_67c367cd (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[75]),
    .e(al_3e0d53ab[91]),
    .f(al_3e0d53ab[123]),
    .o(al_f679ae98));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_1999fd69 (
    .a(al_f679ae98),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[91]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_8a876f90 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[76]),
    .e(al_3e0d53ab[92]),
    .f(al_3e0d53ab[124]),
    .o(al_54c46837));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_16120988 (
    .a(al_54c46837),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[92]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_b4246b20 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[77]),
    .e(al_3e0d53ab[93]),
    .f(al_3e0d53ab[125]),
    .o(al_f6c5d1c0));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6cf54611 (
    .a(al_f6c5d1c0),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[93]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_8fc80e68 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[78]),
    .e(al_3e0d53ab[94]),
    .f(al_3e0d53ab[126]),
    .o(al_70d8d4e8));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_87b9de1b (
    .a(al_70d8d4e8),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[94]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_7cb80a2f (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[79]),
    .e(al_3e0d53ab[95]),
    .f(al_3e0d53ab[127]),
    .o(al_dd59d44c));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_eedc5255 (
    .a(al_dd59d44c),
    .b(al_1f7c5f81),
    .o(al_2982a0b8[95]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_a46ec1eb (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[80]),
    .e(al_3e0d53ab[96]),
    .o(al_2982a0b8[96]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_77f48570 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[81]),
    .e(al_3e0d53ab[97]),
    .o(al_2982a0b8[97]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_b0f3d73 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[82]),
    .e(al_3e0d53ab[98]),
    .o(al_2982a0b8[98]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_f0bf9e6d (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[83]),
    .e(al_3e0d53ab[99]),
    .o(al_2982a0b8[99]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_b8a1bae9 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[148]),
    .e(al_3e0d53ab[164]),
    .o(al_cde313f8[100]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_dc2eb698 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[149]),
    .e(al_3e0d53ab[165]),
    .o(al_cde313f8[101]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c3c96e5f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[150]),
    .e(al_3e0d53ab[166]),
    .o(al_cde313f8[102]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_23a1f26 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[151]),
    .e(al_3e0d53ab[167]),
    .o(al_cde313f8[103]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_66ab43fd (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[152]),
    .e(al_3e0d53ab[168]),
    .o(al_cde313f8[104]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_21a8fea3 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[153]),
    .e(al_3e0d53ab[169]),
    .o(al_cde313f8[105]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_fa9cdfd4 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[154]),
    .e(al_3e0d53ab[170]),
    .o(al_cde313f8[106]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c223ff7d (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[155]),
    .e(al_3e0d53ab[171]),
    .o(al_cde313f8[107]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_eb45a7f6 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[156]),
    .e(al_3e0d53ab[172]),
    .o(al_cde313f8[108]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_7af18319 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[157]),
    .e(al_3e0d53ab[173]),
    .o(al_cde313f8[109]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_a9eabaf6 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[158]),
    .e(al_3e0d53ab[174]),
    .o(al_cde313f8[110]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_33528794 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[159]),
    .e(al_3e0d53ab[175]),
    .o(al_cde313f8[111]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_48d8e37 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[160]),
    .e(al_3e0d53ab[176]),
    .o(al_cde313f8[112]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_ed387634 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[161]),
    .e(al_3e0d53ab[177]),
    .o(al_cde313f8[113]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_7deba3bf (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[162]),
    .e(al_3e0d53ab[178]),
    .o(al_cde313f8[114]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_5af61584 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[163]),
    .e(al_3e0d53ab[179]),
    .o(al_cde313f8[115]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_3176fd6f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[164]),
    .e(al_3e0d53ab[180]),
    .o(al_cde313f8[116]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_e3f8d2e4 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[165]),
    .e(al_3e0d53ab[181]),
    .o(al_cde313f8[117]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_4171cc27 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[166]),
    .e(al_3e0d53ab[182]),
    .o(al_cde313f8[118]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_918bf053 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[167]),
    .e(al_3e0d53ab[183]),
    .o(al_cde313f8[119]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_b3c3dadb (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[168]),
    .e(al_3e0d53ab[184]),
    .o(al_cde313f8[120]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_d7c2ccf4 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[169]),
    .e(al_3e0d53ab[185]),
    .o(al_cde313f8[121]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_f5d1c4e0 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[170]),
    .e(al_3e0d53ab[186]),
    .o(al_cde313f8[122]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_2a54178f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[171]),
    .e(al_3e0d53ab[187]),
    .o(al_cde313f8[123]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_92dd5f68 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[172]),
    .e(al_3e0d53ab[188]),
    .o(al_cde313f8[124]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_ec6f25be (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[173]),
    .e(al_3e0d53ab[189]),
    .o(al_cde313f8[125]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_e480cbfe (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[174]),
    .e(al_3e0d53ab[190]),
    .o(al_cde313f8[126]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_dc4bb525 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[175]),
    .e(al_3e0d53ab[191]),
    .o(al_cde313f8[127]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_eb006bfb (
    .a(al_25e28b94),
    .b(al_e3f231cd[96]),
    .c(al_3e0d53ab[128]),
    .o(al_cde313f8[32]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_76efd1b1 (
    .a(al_25e28b94),
    .b(al_e3f231cd[97]),
    .c(al_3e0d53ab[129]),
    .o(al_cde313f8[33]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_a24d7c03 (
    .a(al_25e28b94),
    .b(al_e3f231cd[98]),
    .c(al_3e0d53ab[130]),
    .o(al_cde313f8[34]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_5becbc7 (
    .a(al_25e28b94),
    .b(al_e3f231cd[99]),
    .c(al_3e0d53ab[131]),
    .o(al_cde313f8[35]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_f51c7863 (
    .a(al_25e28b94),
    .b(al_e3f231cd[100]),
    .c(al_3e0d53ab[132]),
    .o(al_cde313f8[36]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_2f823699 (
    .a(al_25e28b94),
    .b(al_e3f231cd[101]),
    .c(al_3e0d53ab[133]),
    .o(al_cde313f8[37]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_57e4e98a (
    .a(al_25e28b94),
    .b(al_e3f231cd[102]),
    .c(al_3e0d53ab[134]),
    .o(al_cde313f8[38]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_1908f79b (
    .a(al_25e28b94),
    .b(al_e3f231cd[103]),
    .c(al_3e0d53ab[135]),
    .o(al_cde313f8[39]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_901fbff3 (
    .a(al_25e28b94),
    .b(al_e3f231cd[104]),
    .c(al_3e0d53ab[136]),
    .o(al_cde313f8[40]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_2aeaf193 (
    .a(al_25e28b94),
    .b(al_e3f231cd[105]),
    .c(al_3e0d53ab[137]),
    .o(al_cde313f8[41]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_33cd3eb2 (
    .a(al_25e28b94),
    .b(al_e3f231cd[106]),
    .c(al_3e0d53ab[138]),
    .o(al_cde313f8[42]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_2980959c (
    .a(al_25e28b94),
    .b(al_e3f231cd[107]),
    .c(al_3e0d53ab[139]),
    .o(al_cde313f8[43]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9f523492 (
    .a(al_25e28b94),
    .b(al_e3f231cd[108]),
    .c(al_3e0d53ab[140]),
    .o(al_cde313f8[44]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_e6bc26ea (
    .a(al_25e28b94),
    .b(al_e3f231cd[109]),
    .c(al_3e0d53ab[141]),
    .o(al_cde313f8[45]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_ee685ac1 (
    .a(al_25e28b94),
    .b(al_e3f231cd[110]),
    .c(al_3e0d53ab[142]),
    .o(al_cde313f8[46]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_50ac4739 (
    .a(al_25e28b94),
    .b(al_e3f231cd[111]),
    .c(al_3e0d53ab[143]),
    .o(al_cde313f8[47]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9d6776d0 (
    .a(al_25e28b94),
    .b(al_e3f231cd[112]),
    .c(al_3e0d53ab[144]),
    .o(al_cde313f8[48]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_c59b956e (
    .a(al_25e28b94),
    .b(al_e3f231cd[113]),
    .c(al_3e0d53ab[145]),
    .o(al_cde313f8[49]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_84763d3a (
    .a(al_25e28b94),
    .b(al_e3f231cd[114]),
    .c(al_3e0d53ab[146]),
    .o(al_cde313f8[50]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_5d804ef7 (
    .a(al_25e28b94),
    .b(al_e3f231cd[115]),
    .c(al_3e0d53ab[147]),
    .o(al_cde313f8[51]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_47e144b0 (
    .a(al_25e28b94),
    .b(al_e3f231cd[116]),
    .c(al_3e0d53ab[148]),
    .o(al_cde313f8[52]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_dfdd550a (
    .a(al_25e28b94),
    .b(al_e3f231cd[117]),
    .c(al_3e0d53ab[149]),
    .o(al_cde313f8[53]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_6ad6914d (
    .a(al_25e28b94),
    .b(al_e3f231cd[118]),
    .c(al_3e0d53ab[150]),
    .o(al_cde313f8[54]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_e28a92e4 (
    .a(al_25e28b94),
    .b(al_e3f231cd[119]),
    .c(al_3e0d53ab[151]),
    .o(al_cde313f8[55]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_1c124c8c (
    .a(al_25e28b94),
    .b(al_e3f231cd[120]),
    .c(al_3e0d53ab[152]),
    .o(al_cde313f8[56]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_4a2be56a (
    .a(al_25e28b94),
    .b(al_e3f231cd[121]),
    .c(al_3e0d53ab[153]),
    .o(al_cde313f8[57]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_d24cd5d8 (
    .a(al_25e28b94),
    .b(al_e3f231cd[122]),
    .c(al_3e0d53ab[154]),
    .o(al_cde313f8[58]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9f139c22 (
    .a(al_25e28b94),
    .b(al_e3f231cd[123]),
    .c(al_3e0d53ab[155]),
    .o(al_cde313f8[59]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_eee81a89 (
    .a(al_25e28b94),
    .b(al_e3f231cd[124]),
    .c(al_3e0d53ab[156]),
    .o(al_cde313f8[60]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_84ce437 (
    .a(al_25e28b94),
    .b(al_e3f231cd[125]),
    .c(al_3e0d53ab[157]),
    .o(al_cde313f8[61]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_2b821fca (
    .a(al_25e28b94),
    .b(al_e3f231cd[126]),
    .c(al_3e0d53ab[158]),
    .o(al_cde313f8[62]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_c3743771 (
    .a(al_25e28b94),
    .b(al_e3f231cd[127]),
    .c(al_3e0d53ab[159]),
    .o(al_cde313f8[63]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_6dfec8e8 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[128]),
    .e(al_3e0d53ab[160]),
    .o(al_cde313f8[64]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_d1624ed0 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[129]),
    .e(al_3e0d53ab[161]),
    .o(al_cde313f8[65]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_d6a64b63 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[130]),
    .e(al_3e0d53ab[162]),
    .o(al_cde313f8[66]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_ad8ac3e1 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[131]),
    .e(al_3e0d53ab[163]),
    .o(al_cde313f8[67]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_bacc0166 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[132]),
    .e(al_3e0d53ab[164]),
    .o(al_cde313f8[68]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_17a3ef8d (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[133]),
    .e(al_3e0d53ab[165]),
    .o(al_cde313f8[69]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_8d4eed05 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[134]),
    .e(al_3e0d53ab[166]),
    .o(al_cde313f8[70]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_8f89018 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[135]),
    .e(al_3e0d53ab[167]),
    .o(al_cde313f8[71]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_d55f5b07 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[136]),
    .e(al_3e0d53ab[168]),
    .o(al_cde313f8[72]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_af409456 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[137]),
    .e(al_3e0d53ab[169]),
    .o(al_cde313f8[73]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_6c574038 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[138]),
    .e(al_3e0d53ab[170]),
    .o(al_cde313f8[74]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_ba1c7f67 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[139]),
    .e(al_3e0d53ab[171]),
    .o(al_cde313f8[75]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_f3fcb262 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[140]),
    .e(al_3e0d53ab[172]),
    .o(al_cde313f8[76]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_e4e3f4fd (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[141]),
    .e(al_3e0d53ab[173]),
    .o(al_cde313f8[77]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_31ccf485 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[142]),
    .e(al_3e0d53ab[174]),
    .o(al_cde313f8[78]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_9dda6adf (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[143]),
    .e(al_3e0d53ab[175]),
    .o(al_cde313f8[79]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_2c65c31 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[128]),
    .e(al_3e0d53ab[144]),
    .f(al_3e0d53ab[176]),
    .o(al_f59dd527));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_81ad4c95 (
    .a(al_f59dd527),
    .b(al_1f7c5f81),
    .o(al_cde313f8[80]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_477911ed (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[129]),
    .e(al_3e0d53ab[145]),
    .f(al_3e0d53ab[177]),
    .o(al_1975efd7));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_40afe3b (
    .a(al_1975efd7),
    .b(al_1f7c5f81),
    .o(al_cde313f8[81]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_6deeed9e (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[130]),
    .e(al_3e0d53ab[146]),
    .f(al_3e0d53ab[178]),
    .o(al_88804612));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_151db389 (
    .a(al_88804612),
    .b(al_1f7c5f81),
    .o(al_cde313f8[82]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_166da6c (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[131]),
    .e(al_3e0d53ab[147]),
    .f(al_3e0d53ab[179]),
    .o(al_76d4d32b));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_2efb4067 (
    .a(al_76d4d32b),
    .b(al_1f7c5f81),
    .o(al_cde313f8[83]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_8101b067 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[132]),
    .e(al_3e0d53ab[148]),
    .f(al_3e0d53ab[180]),
    .o(al_f748f766));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_90234eb2 (
    .a(al_f748f766),
    .b(al_1f7c5f81),
    .o(al_cde313f8[84]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_cb3786a3 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[133]),
    .e(al_3e0d53ab[149]),
    .f(al_3e0d53ab[181]),
    .o(al_961ce596));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f6ab88eb (
    .a(al_961ce596),
    .b(al_1f7c5f81),
    .o(al_cde313f8[85]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_7022c723 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[134]),
    .e(al_3e0d53ab[150]),
    .f(al_3e0d53ab[182]),
    .o(al_cd1b2b40));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f1d01dd4 (
    .a(al_cd1b2b40),
    .b(al_1f7c5f81),
    .o(al_cde313f8[86]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_662e439a (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[135]),
    .e(al_3e0d53ab[151]),
    .f(al_3e0d53ab[183]),
    .o(al_be7ae2e2));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c61e3768 (
    .a(al_be7ae2e2),
    .b(al_1f7c5f81),
    .o(al_cde313f8[87]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_7f11fb2e (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[136]),
    .e(al_3e0d53ab[152]),
    .f(al_3e0d53ab[184]),
    .o(al_b25b5a5a));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c42c95a6 (
    .a(al_b25b5a5a),
    .b(al_1f7c5f81),
    .o(al_cde313f8[88]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_14ca984f (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[137]),
    .e(al_3e0d53ab[153]),
    .f(al_3e0d53ab[185]),
    .o(al_20384508));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fa2da292 (
    .a(al_20384508),
    .b(al_1f7c5f81),
    .o(al_cde313f8[89]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_3df54b9a (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[138]),
    .e(al_3e0d53ab[154]),
    .f(al_3e0d53ab[186]),
    .o(al_f3f27b05));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_a6f6d20f (
    .a(al_f3f27b05),
    .b(al_1f7c5f81),
    .o(al_cde313f8[90]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_b45900e4 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[139]),
    .e(al_3e0d53ab[155]),
    .f(al_3e0d53ab[187]),
    .o(al_9bc80d94));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b03d2f1c (
    .a(al_9bc80d94),
    .b(al_1f7c5f81),
    .o(al_cde313f8[91]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_961ad455 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[140]),
    .e(al_3e0d53ab[156]),
    .f(al_3e0d53ab[188]),
    .o(al_bb6e492e));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_2e9cef6b (
    .a(al_bb6e492e),
    .b(al_1f7c5f81),
    .o(al_cde313f8[92]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_f146f5f4 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[141]),
    .e(al_3e0d53ab[157]),
    .f(al_3e0d53ab[189]),
    .o(al_867a962f));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_53ed6c31 (
    .a(al_867a962f),
    .b(al_1f7c5f81),
    .o(al_cde313f8[93]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_d0526893 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[142]),
    .e(al_3e0d53ab[158]),
    .f(al_3e0d53ab[190]),
    .o(al_23bdcd5d));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e4f19d24 (
    .a(al_23bdcd5d),
    .b(al_1f7c5f81),
    .o(al_cde313f8[94]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_48a9e8e7 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[143]),
    .e(al_3e0d53ab[159]),
    .f(al_3e0d53ab[191]),
    .o(al_5c5f6698));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_af6ee51a (
    .a(al_5c5f6698),
    .b(al_1f7c5f81),
    .o(al_cde313f8[95]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_d8696111 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[144]),
    .e(al_3e0d53ab[160]),
    .o(al_cde313f8[96]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_f170c8b5 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[145]),
    .e(al_3e0d53ab[161]),
    .o(al_cde313f8[97]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_e5940059 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[146]),
    .e(al_3e0d53ab[162]),
    .o(al_cde313f8[98]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_8a118c68 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[147]),
    .e(al_3e0d53ab[163]),
    .o(al_cde313f8[99]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_6a9fee5c (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[212]),
    .e(al_3e0d53ab[228]),
    .o(al_b43737f6[100]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_cc447f18 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[213]),
    .e(al_3e0d53ab[229]),
    .o(al_b43737f6[101]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c2554202 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[214]),
    .e(al_3e0d53ab[230]),
    .o(al_b43737f6[102]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_28718059 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[215]),
    .e(al_3e0d53ab[231]),
    .o(al_b43737f6[103]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c7f94f9 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[216]),
    .e(al_3e0d53ab[232]),
    .o(al_b43737f6[104]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_aaca9d77 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[217]),
    .e(al_3e0d53ab[233]),
    .o(al_b43737f6[105]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_42a4690d (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[218]),
    .e(al_3e0d53ab[234]),
    .o(al_b43737f6[106]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_f8372972 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[219]),
    .e(al_3e0d53ab[235]),
    .o(al_b43737f6[107]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_9f56d350 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[220]),
    .e(al_3e0d53ab[236]),
    .o(al_b43737f6[108]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_673144e1 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[221]),
    .e(al_3e0d53ab[237]),
    .o(al_b43737f6[109]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_987d2f3a (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[222]),
    .e(al_3e0d53ab[238]),
    .o(al_b43737f6[110]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_8682f165 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[223]),
    .e(al_3e0d53ab[239]),
    .o(al_b43737f6[111]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_3ef87af0 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[224]),
    .e(al_3e0d53ab[240]),
    .o(al_b43737f6[112]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_ab62f5e4 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[225]),
    .e(al_3e0d53ab[241]),
    .o(al_b43737f6[113]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_3cfc9ee3 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[226]),
    .e(al_3e0d53ab[242]),
    .o(al_b43737f6[114]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_a3ae7e92 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[227]),
    .e(al_3e0d53ab[243]),
    .o(al_b43737f6[115]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_3838babd (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[228]),
    .e(al_3e0d53ab[244]),
    .o(al_b43737f6[116]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_75f9c2e7 (
    .a(al_1fba6212),
    .b(al_1f7c5f81),
    .o(al_3c7d7d5c));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_be4dec29 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[229]),
    .e(al_3e0d53ab[245]),
    .o(al_b43737f6[117]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_90cac95f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[230]),
    .e(al_3e0d53ab[246]),
    .o(al_b43737f6[118]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_e706762f (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[231]),
    .e(al_3e0d53ab[247]),
    .o(al_b43737f6[119]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_362688cc (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[232]),
    .e(al_3e0d53ab[248]),
    .o(al_b43737f6[120]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_a46f2cbb (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[233]),
    .e(al_3e0d53ab[249]),
    .o(al_b43737f6[121]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_7d91cfad (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[234]),
    .e(al_3e0d53ab[250]),
    .o(al_b43737f6[122]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_eec4f3eb (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[235]),
    .e(al_3e0d53ab[251]),
    .o(al_b43737f6[123]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_313839c1 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[236]),
    .e(al_3e0d53ab[252]),
    .o(al_b43737f6[124]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_ab9986e1 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[237]),
    .e(al_3e0d53ab[253]),
    .o(al_b43737f6[125]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_334dd162 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[238]),
    .e(al_3e0d53ab[254]),
    .o(al_b43737f6[126]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c989d4cf (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[239]),
    .e(al_3e0d53ab[255]),
    .o(al_b43737f6[127]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_57405135 (
    .a(al_25e28b94),
    .b(al_a1c5f121[96]),
    .c(al_3e0d53ab[192]),
    .o(al_b43737f6[32]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_c6f771d8 (
    .a(al_25e28b94),
    .b(al_a1c5f121[97]),
    .c(al_3e0d53ab[193]),
    .o(al_b43737f6[33]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_e2eb6561 (
    .a(al_25e28b94),
    .b(al_a1c5f121[98]),
    .c(al_3e0d53ab[194]),
    .o(al_b43737f6[34]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_decc31a3 (
    .a(al_25e28b94),
    .b(al_a1c5f121[99]),
    .c(al_3e0d53ab[195]),
    .o(al_b43737f6[35]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_ec14a991 (
    .a(al_25e28b94),
    .b(al_a1c5f121[100]),
    .c(al_3e0d53ab[196]),
    .o(al_b43737f6[36]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_358aff9d (
    .a(al_25e28b94),
    .b(al_a1c5f121[101]),
    .c(al_3e0d53ab[197]),
    .o(al_b43737f6[37]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_7375b8c4 (
    .a(al_25e28b94),
    .b(al_a1c5f121[102]),
    .c(al_3e0d53ab[198]),
    .o(al_b43737f6[38]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9d5df9dc (
    .a(al_25e28b94),
    .b(al_a1c5f121[103]),
    .c(al_3e0d53ab[199]),
    .o(al_b43737f6[39]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_2e4b608a (
    .a(al_25e28b94),
    .b(al_a1c5f121[104]),
    .c(al_3e0d53ab[200]),
    .o(al_b43737f6[40]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_b47df720 (
    .a(al_25e28b94),
    .b(al_a1c5f121[105]),
    .c(al_3e0d53ab[201]),
    .o(al_b43737f6[41]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_edf2a440 (
    .a(al_25e28b94),
    .b(al_a1c5f121[106]),
    .c(al_3e0d53ab[202]),
    .o(al_b43737f6[42]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_7494258d (
    .a(al_25e28b94),
    .b(al_a1c5f121[107]),
    .c(al_3e0d53ab[203]),
    .o(al_b43737f6[43]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_480560fb (
    .a(al_25e28b94),
    .b(al_a1c5f121[108]),
    .c(al_3e0d53ab[204]),
    .o(al_b43737f6[44]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_5cba82e6 (
    .a(al_25e28b94),
    .b(al_a1c5f121[109]),
    .c(al_3e0d53ab[205]),
    .o(al_b43737f6[45]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_a3ed1d15 (
    .a(al_25e28b94),
    .b(al_a1c5f121[110]),
    .c(al_3e0d53ab[206]),
    .o(al_b43737f6[46]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9aa0e0cb (
    .a(al_25e28b94),
    .b(al_a1c5f121[111]),
    .c(al_3e0d53ab[207]),
    .o(al_b43737f6[47]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_74761eda (
    .a(al_25e28b94),
    .b(al_a1c5f121[112]),
    .c(al_3e0d53ab[208]),
    .o(al_b43737f6[48]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_494d3442 (
    .a(al_25e28b94),
    .b(al_a1c5f121[113]),
    .c(al_3e0d53ab[209]),
    .o(al_b43737f6[49]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_743ea2f0 (
    .a(al_25e28b94),
    .b(al_a1c5f121[114]),
    .c(al_3e0d53ab[210]),
    .o(al_b43737f6[50]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_a684d605 (
    .a(al_25e28b94),
    .b(al_a1c5f121[115]),
    .c(al_3e0d53ab[211]),
    .o(al_b43737f6[51]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_fffc3e28 (
    .a(al_25e28b94),
    .b(al_a1c5f121[116]),
    .c(al_3e0d53ab[212]),
    .o(al_b43737f6[52]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9f1c7099 (
    .a(al_25e28b94),
    .b(al_a1c5f121[117]),
    .c(al_3e0d53ab[213]),
    .o(al_b43737f6[53]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_1716403d (
    .a(al_25e28b94),
    .b(al_a1c5f121[118]),
    .c(al_3e0d53ab[214]),
    .o(al_b43737f6[54]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_b149a2c9 (
    .a(al_25e28b94),
    .b(al_a1c5f121[119]),
    .c(al_3e0d53ab[215]),
    .o(al_b43737f6[55]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_c6f0f59 (
    .a(al_25e28b94),
    .b(al_a1c5f121[120]),
    .c(al_3e0d53ab[216]),
    .o(al_b43737f6[56]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_33f1de74 (
    .a(al_25e28b94),
    .b(al_a1c5f121[121]),
    .c(al_3e0d53ab[217]),
    .o(al_b43737f6[57]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_ec4cb628 (
    .a(al_25e28b94),
    .b(al_a1c5f121[122]),
    .c(al_3e0d53ab[218]),
    .o(al_b43737f6[58]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_99060afb (
    .a(al_25e28b94),
    .b(al_a1c5f121[123]),
    .c(al_3e0d53ab[219]),
    .o(al_b43737f6[59]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_1d5c331a (
    .a(al_25e28b94),
    .b(al_a1c5f121[124]),
    .c(al_3e0d53ab[220]),
    .o(al_b43737f6[60]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_3cde6846 (
    .a(al_25e28b94),
    .b(al_a1c5f121[125]),
    .c(al_3e0d53ab[221]),
    .o(al_b43737f6[61]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_2d97487 (
    .a(al_25e28b94),
    .b(al_a1c5f121[126]),
    .c(al_3e0d53ab[222]),
    .o(al_b43737f6[62]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_8addd30d (
    .a(al_25e28b94),
    .b(al_a1c5f121[127]),
    .c(al_3e0d53ab[223]),
    .o(al_b43737f6[63]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_f5c028f5 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[192]),
    .e(al_3e0d53ab[224]),
    .o(al_b43737f6[64]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_1142236f (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[193]),
    .e(al_3e0d53ab[225]),
    .o(al_b43737f6[65]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_746af79 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[194]),
    .e(al_3e0d53ab[226]),
    .o(al_b43737f6[66]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_a3f69a6a (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[195]),
    .e(al_3e0d53ab[227]),
    .o(al_b43737f6[67]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_2b4175de (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[196]),
    .e(al_3e0d53ab[228]),
    .o(al_b43737f6[68]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_59ae85ba (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[197]),
    .e(al_3e0d53ab[229]),
    .o(al_b43737f6[69]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_25b3ae7f (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[198]),
    .e(al_3e0d53ab[230]),
    .o(al_b43737f6[70]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_3a72dabc (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[199]),
    .e(al_3e0d53ab[231]),
    .o(al_b43737f6[71]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_1c2a86a1 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[200]),
    .e(al_3e0d53ab[232]),
    .o(al_b43737f6[72]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_1572ba14 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[201]),
    .e(al_3e0d53ab[233]),
    .o(al_b43737f6[73]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_f334dd45 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[202]),
    .e(al_3e0d53ab[234]),
    .o(al_b43737f6[74]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_49514aec (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[203]),
    .e(al_3e0d53ab[235]),
    .o(al_b43737f6[75]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_2d5d234a (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[204]),
    .e(al_3e0d53ab[236]),
    .o(al_b43737f6[76]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_f3911df0 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[205]),
    .e(al_3e0d53ab[237]),
    .o(al_b43737f6[77]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_ee0cb94f (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[206]),
    .e(al_3e0d53ab[238]),
    .o(al_b43737f6[78]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_9d9ef775 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[207]),
    .e(al_3e0d53ab[239]),
    .o(al_b43737f6[79]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_bc212671 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[192]),
    .e(al_3e0d53ab[208]),
    .f(al_3e0d53ab[240]),
    .o(al_4a2d2508));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_707ff5bf (
    .a(al_4a2d2508),
    .b(al_1f7c5f81),
    .o(al_b43737f6[80]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_f6c1beba (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[193]),
    .e(al_3e0d53ab[209]),
    .f(al_3e0d53ab[241]),
    .o(al_8b27a255));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_bd89d33b (
    .a(al_8b27a255),
    .b(al_1f7c5f81),
    .o(al_b43737f6[81]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_9dd8962c (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[194]),
    .e(al_3e0d53ab[210]),
    .f(al_3e0d53ab[242]),
    .o(al_d31ef303));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_a5b52547 (
    .a(al_d31ef303),
    .b(al_1f7c5f81),
    .o(al_b43737f6[82]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_6cbf7a1f (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[195]),
    .e(al_3e0d53ab[211]),
    .f(al_3e0d53ab[243]),
    .o(al_8d596be2));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3b4c8869 (
    .a(al_8d596be2),
    .b(al_1f7c5f81),
    .o(al_b43737f6[83]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_cff4b0ae (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[196]),
    .e(al_3e0d53ab[212]),
    .f(al_3e0d53ab[244]),
    .o(al_5acc3a2f));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b775b95d (
    .a(al_5acc3a2f),
    .b(al_1f7c5f81),
    .o(al_b43737f6[84]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_7e96862 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[197]),
    .e(al_3e0d53ab[213]),
    .f(al_3e0d53ab[245]),
    .o(al_2244f12b));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_16583c10 (
    .a(al_2244f12b),
    .b(al_1f7c5f81),
    .o(al_b43737f6[85]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_a6c75fbd (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[198]),
    .e(al_3e0d53ab[214]),
    .f(al_3e0d53ab[246]),
    .o(al_ce58a1e1));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_804249c7 (
    .a(al_ce58a1e1),
    .b(al_1f7c5f81),
    .o(al_b43737f6[86]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_d6204993 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[199]),
    .e(al_3e0d53ab[215]),
    .f(al_3e0d53ab[247]),
    .o(al_aa2163c2));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c0c104c1 (
    .a(al_aa2163c2),
    .b(al_1f7c5f81),
    .o(al_b43737f6[87]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_e9dd59f7 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[200]),
    .e(al_3e0d53ab[216]),
    .f(al_3e0d53ab[248]),
    .o(al_42b48cc4));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_a03ebdc1 (
    .a(al_42b48cc4),
    .b(al_1f7c5f81),
    .o(al_b43737f6[88]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_f39c0fc8 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[201]),
    .e(al_3e0d53ab[217]),
    .f(al_3e0d53ab[249]),
    .o(al_4463b457));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_4f26cbcf (
    .a(al_4463b457),
    .b(al_1f7c5f81),
    .o(al_b43737f6[89]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_a8bee2e3 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[202]),
    .e(al_3e0d53ab[218]),
    .f(al_3e0d53ab[250]),
    .o(al_fad9ab0e));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6372ac48 (
    .a(al_fad9ab0e),
    .b(al_1f7c5f81),
    .o(al_b43737f6[90]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_4f8dc662 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[203]),
    .e(al_3e0d53ab[219]),
    .f(al_3e0d53ab[251]),
    .o(al_a3a81a88));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_669ef1d4 (
    .a(al_a3a81a88),
    .b(al_1f7c5f81),
    .o(al_b43737f6[91]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_25d15fcc (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[204]),
    .e(al_3e0d53ab[220]),
    .f(al_3e0d53ab[252]),
    .o(al_fe36a6e2));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3c46e053 (
    .a(al_fe36a6e2),
    .b(al_1f7c5f81),
    .o(al_b43737f6[92]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_4aadc133 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[205]),
    .e(al_3e0d53ab[221]),
    .f(al_3e0d53ab[253]),
    .o(al_acf97feb));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d4415ef8 (
    .a(al_acf97feb),
    .b(al_1f7c5f81),
    .o(al_b43737f6[93]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_47d42355 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[206]),
    .e(al_3e0d53ab[222]),
    .f(al_3e0d53ab[254]),
    .o(al_548ecc42));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_97864b02 (
    .a(al_548ecc42),
    .b(al_1f7c5f81),
    .o(al_b43737f6[94]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_2c9ea13f (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[207]),
    .e(al_3e0d53ab[223]),
    .f(al_3e0d53ab[255]),
    .o(al_dc53c2f4));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_7265e538 (
    .a(al_dc53c2f4),
    .b(al_1f7c5f81),
    .o(al_b43737f6[95]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_af364511 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[208]),
    .e(al_3e0d53ab[224]),
    .o(al_b43737f6[96]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c077aa7a (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[209]),
    .e(al_3e0d53ab[225]),
    .o(al_b43737f6[97]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_fb5eecf6 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[210]),
    .e(al_3e0d53ab[226]),
    .o(al_b43737f6[98]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_75be77b6 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[211]),
    .e(al_3e0d53ab[227]),
    .o(al_b43737f6[99]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_89391f4 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[20]),
    .e(al_3e0d53ab[36]),
    .o(al_880499db[100]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_9a7642e5 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[21]),
    .e(al_3e0d53ab[37]),
    .o(al_880499db[101]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_542bfc2e (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[22]),
    .e(al_3e0d53ab[38]),
    .o(al_880499db[102]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_84579f6e (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[23]),
    .e(al_3e0d53ab[39]),
    .o(al_880499db[103]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_40835e62 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[24]),
    .e(al_3e0d53ab[40]),
    .o(al_880499db[104]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_9fc4fe7c (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[25]),
    .e(al_3e0d53ab[41]),
    .o(al_880499db[105]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_96771c48 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[26]),
    .e(al_3e0d53ab[42]),
    .o(al_880499db[106]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_7476ffd3 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[27]),
    .e(al_3e0d53ab[43]),
    .o(al_880499db[107]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_858f7942 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[28]),
    .e(al_3e0d53ab[44]),
    .o(al_880499db[108]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_bf901e1 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[29]),
    .e(al_3e0d53ab[45]),
    .o(al_880499db[109]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_ea82cbb9 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[30]),
    .e(al_3e0d53ab[46]),
    .o(al_880499db[110]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_5dfc8024 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[31]),
    .e(al_3e0d53ab[47]),
    .o(al_880499db[111]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_34200327 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[32]),
    .e(al_3e0d53ab[48]),
    .o(al_880499db[112]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_d66655f9 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[33]),
    .e(al_3e0d53ab[49]),
    .o(al_880499db[113]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_a95c830 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[34]),
    .e(al_3e0d53ab[50]),
    .o(al_880499db[114]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_d38400e (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[35]),
    .e(al_3e0d53ab[51]),
    .o(al_880499db[115]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_20f8c248 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[36]),
    .e(al_3e0d53ab[52]),
    .o(al_880499db[116]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_692560e5 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[37]),
    .e(al_3e0d53ab[53]),
    .o(al_880499db[117]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_1a9774d1 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[38]),
    .e(al_3e0d53ab[54]),
    .o(al_880499db[118]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_569399d7 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[39]),
    .e(al_3e0d53ab[55]),
    .o(al_880499db[119]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_155875a9 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[40]),
    .e(al_3e0d53ab[56]),
    .o(al_880499db[120]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_adaa404 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[41]),
    .e(al_3e0d53ab[57]),
    .o(al_880499db[121]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_2890e4e8 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[42]),
    .e(al_3e0d53ab[58]),
    .o(al_880499db[122]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_54ab3a3d (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[43]),
    .e(al_3e0d53ab[59]),
    .o(al_880499db[123]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_8378ff43 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[44]),
    .e(al_3e0d53ab[60]),
    .o(al_880499db[124]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_75c9e838 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[45]),
    .e(al_3e0d53ab[61]),
    .o(al_880499db[125]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_57582649 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[46]),
    .e(al_3e0d53ab[62]),
    .o(al_880499db[126]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_800aa2c (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[47]),
    .e(al_3e0d53ab[63]),
    .o(al_880499db[127]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_3b02f597 (
    .a(al_25e28b94),
    .b(al_32e78cf2[96]),
    .c(al_3e0d53ab[0]),
    .o(al_880499db[32]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_7940c441 (
    .a(al_25e28b94),
    .b(al_32e78cf2[97]),
    .c(al_3e0d53ab[1]),
    .o(al_880499db[33]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_cb985a29 (
    .a(al_25e28b94),
    .b(al_32e78cf2[98]),
    .c(al_3e0d53ab[2]),
    .o(al_880499db[34]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_444b0c75 (
    .a(al_25e28b94),
    .b(al_32e78cf2[99]),
    .c(al_3e0d53ab[3]),
    .o(al_880499db[35]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_638e5f76 (
    .a(al_25e28b94),
    .b(al_32e78cf2[100]),
    .c(al_3e0d53ab[4]),
    .o(al_880499db[36]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_b5b00472 (
    .a(al_25e28b94),
    .b(al_32e78cf2[101]),
    .c(al_3e0d53ab[5]),
    .o(al_880499db[37]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_e30caf11 (
    .a(al_25e28b94),
    .b(al_32e78cf2[102]),
    .c(al_3e0d53ab[6]),
    .o(al_880499db[38]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_926f962a (
    .a(al_25e28b94),
    .b(al_32e78cf2[103]),
    .c(al_3e0d53ab[7]),
    .o(al_880499db[39]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_ecdeff97 (
    .a(al_25e28b94),
    .b(al_32e78cf2[104]),
    .c(al_3e0d53ab[8]),
    .o(al_880499db[40]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_4c3ddfd7 (
    .a(al_25e28b94),
    .b(al_32e78cf2[105]),
    .c(al_3e0d53ab[9]),
    .o(al_880499db[41]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_1f81694a (
    .a(al_25e28b94),
    .b(al_32e78cf2[106]),
    .c(al_3e0d53ab[10]),
    .o(al_880499db[42]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_6a4d3108 (
    .a(al_25e28b94),
    .b(al_32e78cf2[107]),
    .c(al_3e0d53ab[11]),
    .o(al_880499db[43]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_1abcf110 (
    .a(al_25e28b94),
    .b(al_32e78cf2[108]),
    .c(al_3e0d53ab[12]),
    .o(al_880499db[44]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_fd0d16f4 (
    .a(al_25e28b94),
    .b(al_32e78cf2[109]),
    .c(al_3e0d53ab[13]),
    .o(al_880499db[45]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_55789fae (
    .a(al_25e28b94),
    .b(al_32e78cf2[110]),
    .c(al_3e0d53ab[14]),
    .o(al_880499db[46]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_88c5660d (
    .a(al_25e28b94),
    .b(al_32e78cf2[111]),
    .c(al_3e0d53ab[15]),
    .o(al_880499db[47]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_4c4966e (
    .a(al_25e28b94),
    .b(al_32e78cf2[112]),
    .c(al_3e0d53ab[16]),
    .o(al_880499db[48]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_2d3080dc (
    .a(al_25e28b94),
    .b(al_32e78cf2[113]),
    .c(al_3e0d53ab[17]),
    .o(al_880499db[49]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_cfaa2a00 (
    .a(al_25e28b94),
    .b(al_32e78cf2[114]),
    .c(al_3e0d53ab[18]),
    .o(al_880499db[50]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_3582d480 (
    .a(al_25e28b94),
    .b(al_32e78cf2[115]),
    .c(al_3e0d53ab[19]),
    .o(al_880499db[51]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_6c962034 (
    .a(al_25e28b94),
    .b(al_32e78cf2[116]),
    .c(al_3e0d53ab[20]),
    .o(al_880499db[52]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_55f3aa8c (
    .a(al_25e28b94),
    .b(al_32e78cf2[117]),
    .c(al_3e0d53ab[21]),
    .o(al_880499db[53]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_30760bf8 (
    .a(al_25e28b94),
    .b(al_32e78cf2[118]),
    .c(al_3e0d53ab[22]),
    .o(al_880499db[54]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_35e9becb (
    .a(al_25e28b94),
    .b(al_32e78cf2[119]),
    .c(al_3e0d53ab[23]),
    .o(al_880499db[55]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_b7d0a8cb (
    .a(al_25e28b94),
    .b(al_32e78cf2[120]),
    .c(al_3e0d53ab[24]),
    .o(al_880499db[56]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_60a4ebe5 (
    .a(al_25e28b94),
    .b(al_32e78cf2[121]),
    .c(al_3e0d53ab[25]),
    .o(al_880499db[57]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_b185e86e (
    .a(al_25e28b94),
    .b(al_32e78cf2[122]),
    .c(al_3e0d53ab[26]),
    .o(al_880499db[58]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_be54b1d4 (
    .a(al_25e28b94),
    .b(al_32e78cf2[123]),
    .c(al_3e0d53ab[27]),
    .o(al_880499db[59]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_89aba3f5 (
    .a(al_25e28b94),
    .b(al_32e78cf2[124]),
    .c(al_3e0d53ab[28]),
    .o(al_880499db[60]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_a75f2de0 (
    .a(al_25e28b94),
    .b(al_32e78cf2[125]),
    .c(al_3e0d53ab[29]),
    .o(al_880499db[61]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_2174e9a1 (
    .a(al_25e28b94),
    .b(al_32e78cf2[126]),
    .c(al_3e0d53ab[30]),
    .o(al_880499db[62]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_ea9371b6 (
    .a(al_25e28b94),
    .b(al_32e78cf2[127]),
    .c(al_3e0d53ab[31]),
    .o(al_880499db[63]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_5c67faee (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[0]),
    .e(al_3e0d53ab[32]),
    .o(al_880499db[64]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_2cf21d28 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[1]),
    .e(al_3e0d53ab[33]),
    .o(al_880499db[65]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_92060bbc (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[2]),
    .e(al_3e0d53ab[34]),
    .o(al_880499db[66]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_f439bba9 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[3]),
    .e(al_3e0d53ab[35]),
    .o(al_880499db[67]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_8856ef46 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[4]),
    .e(al_3e0d53ab[36]),
    .o(al_880499db[68]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_93b7ff43 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[5]),
    .e(al_3e0d53ab[37]),
    .o(al_880499db[69]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_16ba2e48 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[6]),
    .e(al_3e0d53ab[38]),
    .o(al_880499db[70]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_bc5d4a50 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[7]),
    .e(al_3e0d53ab[39]),
    .o(al_880499db[71]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_532f186e (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[8]),
    .e(al_3e0d53ab[40]),
    .o(al_880499db[72]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_e0e4078a (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[9]),
    .e(al_3e0d53ab[41]),
    .o(al_880499db[73]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_ed523bd0 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[10]),
    .e(al_3e0d53ab[42]),
    .o(al_880499db[74]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_7daf3947 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[11]),
    .e(al_3e0d53ab[43]),
    .o(al_880499db[75]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_2e96cad6 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[12]),
    .e(al_3e0d53ab[44]),
    .o(al_880499db[76]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_2cfba262 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[13]),
    .e(al_3e0d53ab[45]),
    .o(al_880499db[77]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_cdf3e585 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[14]),
    .e(al_3e0d53ab[46]),
    .o(al_880499db[78]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_9806459d (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[15]),
    .e(al_3e0d53ab[47]),
    .o(al_880499db[79]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_f220ce8a (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[0]),
    .e(al_3e0d53ab[16]),
    .f(al_3e0d53ab[48]),
    .o(al_369dae91));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f027244e (
    .a(al_369dae91),
    .b(al_1f7c5f81),
    .o(al_880499db[80]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_800eced7 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[1]),
    .e(al_3e0d53ab[17]),
    .f(al_3e0d53ab[49]),
    .o(al_fa0877ed));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6733937c (
    .a(al_fa0877ed),
    .b(al_1f7c5f81),
    .o(al_880499db[81]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_e66c21d0 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[2]),
    .e(al_3e0d53ab[18]),
    .f(al_3e0d53ab[50]),
    .o(al_e1e4e320));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3e21d3ad (
    .a(al_e1e4e320),
    .b(al_1f7c5f81),
    .o(al_880499db[82]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_d323af20 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[3]),
    .e(al_3e0d53ab[19]),
    .f(al_3e0d53ab[51]),
    .o(al_d84d421));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ccbf5efc (
    .a(al_d84d421),
    .b(al_1f7c5f81),
    .o(al_880499db[83]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_e68e7b21 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[4]),
    .e(al_3e0d53ab[20]),
    .f(al_3e0d53ab[52]),
    .o(al_12e89d71));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_337ab4be (
    .a(al_12e89d71),
    .b(al_1f7c5f81),
    .o(al_880499db[84]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_7bfab608 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[5]),
    .e(al_3e0d53ab[21]),
    .f(al_3e0d53ab[53]),
    .o(al_a73e260c));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_90905f6b (
    .a(al_a73e260c),
    .b(al_1f7c5f81),
    .o(al_880499db[85]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_b266cd2 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[6]),
    .e(al_3e0d53ab[22]),
    .f(al_3e0d53ab[54]),
    .o(al_b7c175ec));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f106f366 (
    .a(al_b7c175ec),
    .b(al_1f7c5f81),
    .o(al_880499db[86]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_234022e5 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[7]),
    .e(al_3e0d53ab[23]),
    .f(al_3e0d53ab[55]),
    .o(al_a8c83515));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_240829c6 (
    .a(al_a8c83515),
    .b(al_1f7c5f81),
    .o(al_880499db[87]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_29cd8dfe (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[8]),
    .e(al_3e0d53ab[24]),
    .f(al_3e0d53ab[56]),
    .o(al_698080d7));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_80cb283c (
    .a(al_698080d7),
    .b(al_1f7c5f81),
    .o(al_880499db[88]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_59835d5e (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[9]),
    .e(al_3e0d53ab[25]),
    .f(al_3e0d53ab[57]),
    .o(al_ebc69845));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cb24b64d (
    .a(al_ebc69845),
    .b(al_1f7c5f81),
    .o(al_880499db[89]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_8909790e (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[10]),
    .e(al_3e0d53ab[26]),
    .f(al_3e0d53ab[58]),
    .o(al_5949896a));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c8bff187 (
    .a(al_5949896a),
    .b(al_1f7c5f81),
    .o(al_880499db[90]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_c697727c (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[11]),
    .e(al_3e0d53ab[27]),
    .f(al_3e0d53ab[59]),
    .o(al_6ddecd31));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b1b1b06f (
    .a(al_6ddecd31),
    .b(al_1f7c5f81),
    .o(al_880499db[91]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_6ae71fd4 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[12]),
    .e(al_3e0d53ab[28]),
    .f(al_3e0d53ab[60]),
    .o(al_cf8fae09));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_651cfe36 (
    .a(al_cf8fae09),
    .b(al_1f7c5f81),
    .o(al_880499db[92]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_be9b57bc (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[13]),
    .e(al_3e0d53ab[29]),
    .f(al_3e0d53ab[61]),
    .o(al_64c4b1ee));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f1e3a8cb (
    .a(al_64c4b1ee),
    .b(al_1f7c5f81),
    .o(al_880499db[93]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_6a524e8f (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[14]),
    .e(al_3e0d53ab[30]),
    .f(al_3e0d53ab[62]),
    .o(al_1551352));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e01e5a4b (
    .a(al_1551352),
    .b(al_1f7c5f81),
    .o(al_880499db[94]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_6113bc94 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[15]),
    .e(al_3e0d53ab[31]),
    .f(al_3e0d53ab[63]),
    .o(al_2192db1e));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_aaa3708b (
    .a(al_2192db1e),
    .b(al_1f7c5f81),
    .o(al_880499db[95]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_3afc5483 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[16]),
    .e(al_3e0d53ab[32]),
    .o(al_880499db[96]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_afa1d6b2 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[17]),
    .e(al_3e0d53ab[33]),
    .o(al_880499db[97]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_e1276b6c (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[18]),
    .e(al_3e0d53ab[34]),
    .o(al_880499db[98]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_c4638a2e (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[19]),
    .e(al_3e0d53ab[35]),
    .o(al_880499db[99]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~B*~A))"),
    .INIT(16'hff10))
    al_98bd959f (
    .a(al_4732ba15[0]),
    .b(al_4732ba15[1]),
    .c(al_cc4d831c[0]),
    .d(al_8679dfa[8]),
    .o(al_ea19deeb[0]));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*~C*~(~B*~A))"),
    .INIT(64'h00000e0000000000))
    al_c22d649b (
    .a(al_4732ba15[0]),
    .b(al_4732ba15[1]),
    .c(al_72785055[0]),
    .d(al_72785055[2]),
    .e(al_72785055[1]),
    .f(al_cc4d831c[0]),
    .o(al_ea19deeb[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_a5910fd4 (
    .a(al_b4da789e[0]),
    .b(al_b4da789e[1]),
    .o(al_1fba6212));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_d7c72f89 (
    .a(al_d9b4cc10[0]),
    .b(al_d9b4cc10[1]),
    .c(al_d9b4cc10[2]),
    .o(al_4d9c76b0));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_4f667e4e (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[264]),
    .e(al_3e0d53ab[266]),
    .f(al_3e0d53ab[270]),
    .o(al_70c902df));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_93e3215b (
    .a(al_70c902df),
    .b(al_1f7c5f81),
    .o(al_8ef9bc8c[10]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_8d768b6b (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[265]),
    .e(al_3e0d53ab[267]),
    .f(al_3e0d53ab[271]),
    .o(al_56881e67));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_19f87884 (
    .a(al_56881e67),
    .b(al_1f7c5f81),
    .o(al_8ef9bc8c[11]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_552bfcac (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[266]),
    .e(al_3e0d53ab[268]),
    .o(al_8ef9bc8c[12]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_a3dc294d (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[267]),
    .e(al_3e0d53ab[269]),
    .o(al_8ef9bc8c[13]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_b8454ee (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[268]),
    .e(al_3e0d53ab[270]),
    .o(al_8ef9bc8c[14]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_618310f4 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[269]),
    .e(al_3e0d53ab[271]),
    .o(al_8ef9bc8c[15]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_ffd66b3d (
    .a(al_25e28b94),
    .b(al_55ed1bfd[12]),
    .c(al_3e0d53ab[264]),
    .o(al_8ef9bc8c[4]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_502ba324 (
    .a(al_25e28b94),
    .b(al_55ed1bfd[13]),
    .c(al_3e0d53ab[265]),
    .o(al_8ef9bc8c[5]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_c2da2178 (
    .a(al_25e28b94),
    .b(al_55ed1bfd[14]),
    .c(al_3e0d53ab[266]),
    .o(al_8ef9bc8c[6]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_24ba487d (
    .a(al_25e28b94),
    .b(al_55ed1bfd[15]),
    .c(al_3e0d53ab[267]),
    .o(al_8ef9bc8c[7]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_e45b9f30 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[264]),
    .e(al_3e0d53ab[268]),
    .o(al_8ef9bc8c[8]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_dfa41ac6 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[265]),
    .e(al_3e0d53ab[269]),
    .o(al_8ef9bc8c[9]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_ba3478f2 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[272]),
    .e(al_3e0d53ab[274]),
    .f(al_3e0d53ab[278]),
    .o(al_45a1a0f8));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b54f6f94 (
    .a(al_45a1a0f8),
    .b(al_1f7c5f81),
    .o(al_e1aabbd4[10]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_835f64a7 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[273]),
    .e(al_3e0d53ab[275]),
    .f(al_3e0d53ab[279]),
    .o(al_72d2fdcd));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_5fa332ec (
    .a(al_72d2fdcd),
    .b(al_1f7c5f81),
    .o(al_e1aabbd4[11]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_469ef7b1 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[274]),
    .e(al_3e0d53ab[276]),
    .o(al_e1aabbd4[12]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_f07fe7e6 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[275]),
    .e(al_3e0d53ab[277]),
    .o(al_e1aabbd4[13]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_3ba72f7 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[276]),
    .e(al_3e0d53ab[278]),
    .o(al_e1aabbd4[14]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_b1972649 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[277]),
    .e(al_3e0d53ab[279]),
    .o(al_e1aabbd4[15]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_8a03d08d (
    .a(al_25e28b94),
    .b(al_b0d99cb1[12]),
    .c(al_3e0d53ab[272]),
    .o(al_e1aabbd4[4]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_3e32d738 (
    .a(al_25e28b94),
    .b(al_b0d99cb1[13]),
    .c(al_3e0d53ab[273]),
    .o(al_e1aabbd4[5]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_539cd054 (
    .a(al_25e28b94),
    .b(al_b0d99cb1[14]),
    .c(al_3e0d53ab[274]),
    .o(al_e1aabbd4[6]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_a9944580 (
    .a(al_25e28b94),
    .b(al_b0d99cb1[15]),
    .c(al_3e0d53ab[275]),
    .o(al_e1aabbd4[7]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_a1ef55fb (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[272]),
    .e(al_3e0d53ab[276]),
    .o(al_e1aabbd4[8]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_da5be960 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[273]),
    .e(al_3e0d53ab[277]),
    .o(al_e1aabbd4[9]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_1892edc9 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[280]),
    .e(al_3e0d53ab[282]),
    .f(al_3e0d53ab[286]),
    .o(al_45d223ab));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_61054357 (
    .a(al_45d223ab),
    .b(al_1f7c5f81),
    .o(al_4f2a09ff[10]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_7b47bb47 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[281]),
    .e(al_3e0d53ab[283]),
    .f(al_3e0d53ab[287]),
    .o(al_f759090a));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c69128b (
    .a(al_f759090a),
    .b(al_1f7c5f81),
    .o(al_4f2a09ff[11]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_ba8c4f9a (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[282]),
    .e(al_3e0d53ab[284]),
    .o(al_4f2a09ff[12]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_2dbcfca2 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[283]),
    .e(al_3e0d53ab[285]),
    .o(al_4f2a09ff[13]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_53394ee8 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[284]),
    .e(al_3e0d53ab[286]),
    .o(al_4f2a09ff[14]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_3a68c59d (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[285]),
    .e(al_3e0d53ab[287]),
    .o(al_4f2a09ff[15]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_aeb04853 (
    .a(al_25e28b94),
    .b(al_f949a7ee[12]),
    .c(al_3e0d53ab[280]),
    .o(al_4f2a09ff[4]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_6dd359ee (
    .a(al_25e28b94),
    .b(al_f949a7ee[13]),
    .c(al_3e0d53ab[281]),
    .o(al_4f2a09ff[5]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_bf8395b3 (
    .a(al_25e28b94),
    .b(al_f949a7ee[14]),
    .c(al_3e0d53ab[282]),
    .o(al_4f2a09ff[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_a4cf4340 (
    .a(al_1fba6212),
    .b(al_1f7c5f81),
    .o(al_25e28b94));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_eaa4017f (
    .a(al_25e28b94),
    .b(al_f949a7ee[15]),
    .c(al_3e0d53ab[283]),
    .o(al_4f2a09ff[7]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_c15726e8 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[280]),
    .e(al_3e0d53ab[284]),
    .o(al_4f2a09ff[8]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_c90b95f6 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[281]),
    .e(al_3e0d53ab[285]),
    .o(al_4f2a09ff[9]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_e27c7cca (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[256]),
    .e(al_3e0d53ab[258]),
    .f(al_3e0d53ab[262]),
    .o(al_4d6aba82));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_5ce8f937 (
    .a(al_4d6aba82),
    .b(al_1f7c5f81),
    .o(al_523e9f7a[10]));
  AL_MAP_LUT6 #(
    .EQN("~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*~(F)*~(B)+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*~(B)+~((E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C))*F*B+(E*~((D*A))*~(C)+E*(D*A)*~(C)+~(E)*(D*A)*C+E*(D*A)*C)*F*B)"),
    .INIT(64'h10301333dcfcdfff))
    al_d5cf4157 (
    .a(al_4d9c76b0),
    .b(al_1fba6212),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[257]),
    .e(al_3e0d53ab[259]),
    .f(al_3e0d53ab[263]),
    .o(al_790ebcd));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f012aedb (
    .a(al_790ebcd),
    .b(al_1f7c5f81),
    .o(al_523e9f7a[11]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_43f3b1c2 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[258]),
    .e(al_3e0d53ab[260]),
    .o(al_523e9f7a[12]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_34c2b2e9 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[259]),
    .e(al_3e0d53ab[261]),
    .o(al_523e9f7a[13]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_5ac08e12 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[260]),
    .e(al_3e0d53ab[262]),
    .o(al_523e9f7a[14]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E*~((D*B))*~(C)+E*(D*B)*~(C)+~(E)*(D*B)*C+E*(D*B)*C))"),
    .INIT(32'h8a0a8000))
    al_7bb06bb5 (
    .a(al_3c7d7d5c),
    .b(al_4d9c76b0),
    .c(al_48eb6d34[0]),
    .d(al_3e0d53ab[261]),
    .e(al_3e0d53ab[263]),
    .o(al_523e9f7a[15]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_eaa3b819 (
    .a(al_25e28b94),
    .b(al_4340e4e7[12]),
    .c(al_3e0d53ab[256]),
    .o(al_523e9f7a[4]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_6d0c523e (
    .a(al_25e28b94),
    .b(al_4340e4e7[13]),
    .c(al_3e0d53ab[257]),
    .o(al_523e9f7a[5]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_9f5ce277 (
    .a(al_25e28b94),
    .b(al_4340e4e7[14]),
    .c(al_3e0d53ab[258]),
    .o(al_523e9f7a[6]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_1ba5e180 (
    .a(al_25e28b94),
    .b(al_4340e4e7[15]),
    .c(al_3e0d53ab[259]),
    .o(al_523e9f7a[7]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_a5286eb8 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[256]),
    .e(al_3e0d53ab[260]),
    .o(al_523e9f7a[8]));
  AL_MAP_LUT5 #(
    .EQN("(C*((D*~B)*~(E)*~(A)+(D*~B)*E*~(A)+~((D*~B))*E*A+(D*~B)*E*A))"),
    .INIT(32'hb0a01000))
    al_69552a71 (
    .a(al_1fba6212),
    .b(al_48eb6d34[0]),
    .c(al_1f7c5f81),
    .d(al_3e0d53ab[257]),
    .e(al_3e0d53ab[261]),
    .o(al_523e9f7a[9]));
  AL_DFF_0 al_1c750ff1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2ee87d50),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90d84dc7[0]));
  AL_DFF_0 al_d0832055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_91632424),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_71e16f2b));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    al_19410438 (
    .a(al_903070b1),
    .b(init_calib_complete),
    .c(al_90d84dc7[0]),
    .d(al_df80405c),
    .o(al_59addda8));
  AL_MAP_LUT5 #(
    .EQN("(~C*(A*B*~(D)*~(E)+A*B*~(D)*E+~(A)*~(B)*D*E+A*~(B)*D*E))"),
    .INIT(32'h03080008))
    al_a4a39d4d (
    .a(al_aafc78b6),
    .b(al_a67dc86a[0]),
    .c(al_a67dc86a[1]),
    .d(al_a67dc86a[2]),
    .e(al_e620c305),
    .o(al_52665bb8));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    al_b55dff0a (
    .a(al_52665bb8),
    .b(al_71e16f2b),
    .c(al_c360bf4c[0]),
    .o(al_91632424));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_38fef0d7 (
    .a(al_b93da8d5[0]),
    .b(al_b93da8d5[1]),
    .c(al_73f8a8a7[0]),
    .d(al_f0482f12[0]),
    .e(al_f0482f12[1]),
    .o(al_80083fda[0]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_2036a10f (
    .a(al_b93da8d5[0]),
    .b(al_b93da8d5[1]),
    .c(al_73f8a8a7[2]),
    .d(al_a5104c4f[0]),
    .e(al_a5104c4f[1]),
    .o(al_80083fda[2]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_8f28f749 (
    .a(al_b93da8d5[0]),
    .b(al_b93da8d5[1]),
    .c(al_73f8a8a7[1]),
    .d(al_4b620bb0[0]),
    .e(al_4b620bb0[1]),
    .o(al_80083fda[1]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(D*~(F@C)*~(E@B)))"),
    .INIT(64'h1555455551555455))
    al_c4a6229d (
    .a(al_80083fda[2]),
    .b(al_b93da8d5[0]),
    .c(al_b93da8d5[1]),
    .d(al_73f8a8a7[3]),
    .e(al_dac85437[0]),
    .f(al_dac85437[1]),
    .o(al_7a00688b));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_51a8cf12 (
    .a(al_59addda8),
    .b(al_ac74f6f1),
    .o(al_99c9c113));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_a9916d5a (
    .a(al_99c9c113),
    .b(al_7a00688b),
    .c(al_80083fda[0]),
    .d(al_80083fda[1]),
    .o(al_aafc78b6));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*~A))"),
    .INIT(8'hc9))
    al_82bc68b7 (
    .a(al_cfaa4b74),
    .b(al_1c7e0f23),
    .c(al_2b3c55e4),
    .o(al_5d5ab475[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(~D*~B*~A))"),
    .INIT(16'hf0e1))
    al_61eee6ef (
    .a(al_cfaa4b74),
    .b(al_1c7e0f23),
    .c(al_80cba1f),
    .d(al_2b3c55e4),
    .o(al_5d5ab475[2]));
  AL_MAP_LUT6 #(
    .EQN("(E@(~F*~D*~C*~B*~A))"),
    .INIT(64'hffff0000fffe0001))
    al_fb7720f1 (
    .a(al_cfaa4b74),
    .b(al_1c7e0f23),
    .c(al_80cba1f),
    .d(al_2f87218f),
    .e(al_2d60bf7c),
    .f(al_2b3c55e4),
    .o(al_5d5ab475[4]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_27967175 (
    .a(al_cfaa4b74),
    .b(al_2b3c55e4),
    .o(al_5d5ab475[0]));
  AL_MAP_LUT5 #(
    .EQN("(D@(~E*~C*~B*~A))"),
    .INIT(32'hff00fe01))
    al_c88b6fde (
    .a(al_cfaa4b74),
    .b(al_1c7e0f23),
    .c(al_80cba1f),
    .d(al_2f87218f),
    .e(al_2b3c55e4),
    .o(al_5d5ab475[3]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_29f9e23a (
    .a(al_5d5ab475[3]),
    .b(al_5d5ab475[0]),
    .c(al_1c7e0f23),
    .d(al_80cba1f),
    .e(al_2d60bf7c),
    .o(al_d7619b2[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_1168c5cf (
    .a(al_d7619b2[0]),
    .b(al_2b3c55e4),
    .o(al_d549f91e[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_feee6591 (
    .a(al_c2a06982[0]),
    .b(al_c3bcd0f7[0]),
    .c(al_35348eec[0]),
    .d(al_cd4b89ad[0]),
    .e(al_ffbe21a4[0]),
    .f(al_ffbe21a4[1]),
    .o(al_20b2d1cd[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_83a6f728 (
    .a(al_c2a06982[1]),
    .b(al_c3bcd0f7[1]),
    .c(al_35348eec[1]),
    .d(al_cd4b89ad[1]),
    .e(al_ffbe21a4[0]),
    .f(al_ffbe21a4[1]),
    .o(al_20b2d1cd[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_578232f2 (
    .a(al_c2a06982[2]),
    .b(al_c3bcd0f7[2]),
    .c(al_35348eec[2]),
    .d(al_cd4b89ad[2]),
    .e(al_ffbe21a4[0]),
    .f(al_ffbe21a4[1]),
    .o(al_20b2d1cd[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_4a79253c (
    .a(al_c2a06982[3]),
    .b(al_c3bcd0f7[3]),
    .c(al_35348eec[3]),
    .d(al_cd4b89ad[3]),
    .e(al_ffbe21a4[0]),
    .f(al_ffbe21a4[1]),
    .o(al_20b2d1cd[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_d1197a2f (
    .a(al_c2a06982[4]),
    .b(al_c3bcd0f7[4]),
    .c(al_35348eec[4]),
    .d(al_cd4b89ad[4]),
    .e(al_ffbe21a4[0]),
    .f(al_ffbe21a4[1]),
    .o(al_20b2d1cd[4]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    al_5c7716a1 (
    .a(al_1e3dbb5f),
    .b(al_c46598af[0]),
    .c(al_c46598af[1]),
    .o(al_cebaaa2a));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_2754f502 (
    .a(al_cebaaa2a),
    .b(al_ffbe21a4[0]),
    .o(al_d5c3e265[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*~A))"),
    .INIT(8'hb4))
    al_dab13a79 (
    .a(al_cebaaa2a),
    .b(al_ffbe21a4[0]),
    .c(al_ffbe21a4[1]),
    .o(al_d5c3e265[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C@(B*~A))"),
    .INIT(8'h4b))
    al_5313a501 (
    .a(al_8bee4cd6),
    .b(al_954ec2c7),
    .c(al_99c445b5[0]),
    .o(al_765e8240[0]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B*~A)))"),
    .INIT(16'h4fb0))
    al_b8e1d0f4 (
    .a(al_8bee4cd6),
    .b(al_954ec2c7),
    .c(al_99c445b5[0]),
    .d(al_99c445b5[1]),
    .o(al_765e8240[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_9548ebe2 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_d5c3e265[0]),
    .d(al_d5c3e265[1]),
    .o(al_3b2c2aa));
  AL_DFF_0 al_d6d5cb80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3b2c2aa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a415a42));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(C*~A))"),
    .INIT(16'h639c))
    al_38e73661 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_d5c3e265[0]),
    .d(al_d5c3e265[1]),
    .o(al_b37f6146[1]));
  AL_DFF_0 al_73b0671e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b37f6146[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_891340a1));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_1205fcd6 (
    .a(al_99c445b5[0]),
    .b(al_99c445b5[1]),
    .o(al_10206333[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*~A)))"),
    .INIT(16'h004f))
    al_4c022cfd (
    .a(al_8bee4cd6),
    .b(al_954ec2c7),
    .c(al_10206333[0]),
    .d(al_73f8a8a7[0]),
    .o(al_ba9c6360));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*~B))"),
    .INIT(16'h5554))
    al_ffe4e5d9 (
    .a(al_ba9c6360),
    .b(al_cebaaa2a),
    .c(al_ffbe21a4[0]),
    .d(al_ffbe21a4[1]),
    .o(al_845e0bd1[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_ac364abb (
    .a(al_99c445b5[0]),
    .b(al_99c445b5[1]),
    .o(al_10206333[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*~A)))"),
    .INIT(16'h004f))
    al_79c2ee3a (
    .a(al_8bee4cd6),
    .b(al_954ec2c7),
    .c(al_10206333[1]),
    .d(al_73f8a8a7[1]),
    .o(al_22cfe3fb));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*~B))"),
    .INIT(16'h5545))
    al_b21cc237 (
    .a(al_22cfe3fb),
    .b(al_cebaaa2a),
    .c(al_ffbe21a4[0]),
    .d(al_ffbe21a4[1]),
    .o(al_845e0bd1[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3ab0b079 (
    .a(al_99c445b5[0]),
    .b(al_99c445b5[1]),
    .o(al_10206333[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*~A)))"),
    .INIT(16'h004f))
    al_f88f2d10 (
    .a(al_8bee4cd6),
    .b(al_954ec2c7),
    .c(al_10206333[2]),
    .d(al_73f8a8a7[2]),
    .o(al_1f5636ed));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    al_ecc39403 (
    .a(al_1f5636ed),
    .b(al_cebaaa2a),
    .c(al_ffbe21a4[0]),
    .d(al_ffbe21a4[1]),
    .o(al_845e0bd1[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_4dfa615e (
    .a(al_99c445b5[0]),
    .b(al_99c445b5[1]),
    .o(al_10206333[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*~A)))"),
    .INIT(16'h004f))
    al_62a32638 (
    .a(al_8bee4cd6),
    .b(al_954ec2c7),
    .c(al_10206333[3]),
    .d(al_73f8a8a7[3]),
    .o(al_d53d23aa));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    al_5ee23c79 (
    .a(al_d53d23aa),
    .b(al_cebaaa2a),
    .c(al_ffbe21a4[0]),
    .d(al_ffbe21a4[1]),
    .o(al_845e0bd1[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_82b1a929 (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[11]),
    .d(al_4b620bb0[11]),
    .e(al_a5104c4f[11]),
    .f(al_dac85437[11]),
    .o(al_b909a17b));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_dee75a95 (
    .a(al_b909a17b),
    .b(al_8a415a42),
    .c(al_b93da8d5[11]),
    .o(al_71f78ff1[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_366e7201 (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[12]),
    .d(al_4b620bb0[12]),
    .e(al_a5104c4f[12]),
    .f(al_dac85437[12]),
    .o(al_d4376192));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_c132078a (
    .a(al_d4376192),
    .b(al_8a415a42),
    .c(al_b93da8d5[12]),
    .o(al_71f78ff1[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_23f446c3 (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[13]),
    .d(al_4b620bb0[13]),
    .e(al_a5104c4f[13]),
    .f(al_dac85437[13]),
    .o(al_cd1bbfcd));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_e08e0184 (
    .a(al_cd1bbfcd),
    .b(al_8a415a42),
    .c(al_b93da8d5[13]),
    .o(al_71f78ff1[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_6e37bfdc (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[14]),
    .d(al_4b620bb0[14]),
    .e(al_a5104c4f[14]),
    .f(al_dac85437[14]),
    .o(al_45e379c7));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_2dae0f1e (
    .a(al_45e379c7),
    .b(al_8a415a42),
    .c(al_b93da8d5[14]),
    .o(al_71f78ff1[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_492e01e1 (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[15]),
    .d(al_4b620bb0[15]),
    .e(al_a5104c4f[15]),
    .f(al_dac85437[15]),
    .o(al_e4ce0401));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_854385c9 (
    .a(al_e4ce0401),
    .b(al_8a415a42),
    .c(al_b93da8d5[15]),
    .o(al_71f78ff1[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_f65ee865 (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[16]),
    .d(al_4b620bb0[16]),
    .e(al_a5104c4f[16]),
    .f(al_dac85437[16]),
    .o(al_67a5cae3));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_e934f881 (
    .a(al_67a5cae3),
    .b(al_8a415a42),
    .c(al_b93da8d5[16]),
    .o(al_71f78ff1[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_c668398f (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[17]),
    .d(al_4b620bb0[17]),
    .e(al_a5104c4f[17]),
    .f(al_dac85437[17]),
    .o(al_bdd2644));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_801600c2 (
    .a(al_bdd2644),
    .b(al_8a415a42),
    .c(al_b93da8d5[17]),
    .o(al_71f78ff1[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_67749679 (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[2]),
    .d(al_4b620bb0[2]),
    .e(al_a5104c4f[2]),
    .f(al_dac85437[2]),
    .o(al_fc597f88));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_402b0d56 (
    .a(al_fc597f88),
    .b(al_8a415a42),
    .c(al_b93da8d5[2]),
    .o(al_71f78ff1[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_e5ad465 (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[48]),
    .d(al_4b620bb0[48]),
    .e(al_a5104c4f[48]),
    .f(al_dac85437[48]),
    .o(al_7f9b11b5));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_3d03f647 (
    .a(al_7f9b11b5),
    .b(al_8a415a42),
    .c(al_b93da8d5[48]),
    .o(al_71f78ff1[48]));
  AL_DFF_0 al_ca120137 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[48]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_81cbac46[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_5104f56c (
    .a(al_47a64ed5[0]),
    .b(al_75c1ef4c[0]),
    .c(al_ce7d4278[0]),
    .d(al_ad4756a7[0]),
    .e(al_879aba03[0]),
    .f(al_879aba03[1]),
    .o(al_9f407117));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)*~(A)+~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B*~(A)+~(~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*B*A+~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B*A)"),
    .INIT(64'h7777722727722222))
    al_cd5daf2e (
    .a(al_15b16fc6),
    .b(al_9f407117),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[0]),
    .f(al_75c0d27f[0]),
    .o(al_3ee9f2ae[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_4cb05653 (
    .a(al_3ee9f2ae[0]),
    .b(al_75c1ef4c[0]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1f23ce73[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_124aae26 (
    .a(al_3ee9f2ae[0]),
    .b(al_ad4756a7[0]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1bc63bd7[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_2d0edff9 (
    .a(al_3ee9f2ae[0]),
    .b(al_ce7d4278[0]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_abc55d75[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_85b833f2 (
    .a(al_3ee9f2ae[0]),
    .b(al_47a64ed5[0]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_f8f25e7b[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_c37e0ee (
    .a(al_1f23ce73[0]),
    .b(al_1bc63bd7[0]),
    .c(al_abc55d75[0]),
    .d(al_f8f25e7b[0]),
    .e(al_99c445b5[0]),
    .f(al_99c445b5[1]),
    .o(al_b6b411a2[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_f8b38804 (
    .a(al_47a64ed5[1]),
    .b(al_75c1ef4c[1]),
    .c(al_ce7d4278[1]),
    .d(al_ad4756a7[1]),
    .e(al_879aba03[0]),
    .f(al_879aba03[1]),
    .o(al_bfc02a10));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)*~(A)+~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B*~(A)+~(~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*B*A+~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B*A)"),
    .INIT(64'h7777722727722222))
    al_8c9a79e (
    .a(al_15b16fc6),
    .b(al_bfc02a10),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[1]),
    .f(al_75c0d27f[1]),
    .o(al_3ee9f2ae[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_ae03507a (
    .a(al_3ee9f2ae[1]),
    .b(al_75c1ef4c[1]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1f23ce73[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_ef3cdc83 (
    .a(al_3ee9f2ae[1]),
    .b(al_ad4756a7[1]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1bc63bd7[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_b854a180 (
    .a(al_3ee9f2ae[1]),
    .b(al_ce7d4278[1]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_abc55d75[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_d5c23620 (
    .a(al_3ee9f2ae[1]),
    .b(al_47a64ed5[1]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_f8f25e7b[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_8e0e6239 (
    .a(al_1f23ce73[1]),
    .b(al_1bc63bd7[1]),
    .c(al_abc55d75[1]),
    .d(al_f8f25e7b[1]),
    .e(al_99c445b5[0]),
    .f(al_99c445b5[1]),
    .o(al_b6b411a2[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_a97388b2 (
    .a(al_47a64ed5[2]),
    .b(al_75c1ef4c[2]),
    .c(al_ce7d4278[2]),
    .d(al_ad4756a7[2]),
    .e(al_879aba03[0]),
    .f(al_879aba03[1]),
    .o(al_8abd3059));
  AL_MAP_LUT6 #(
    .EQN("(~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)*~(A)+~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B*~(A)+~(~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*B*A+~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B*A)"),
    .INIT(64'h88888dd8d88ddddd))
    al_b9956a62 (
    .a(al_15b16fc6),
    .b(al_8abd3059),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[2]),
    .f(al_75c0d27f[2]),
    .o(al_9b9e072a));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((~D*C))+~B*A*~((~D*C))+~(~B)*A*(~D*C)+~B*A*(~D*C))"),
    .INIT(16'hcc5c))
    al_a95dac84 (
    .a(al_9b9e072a),
    .b(al_75c1ef4c[2]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1f23ce73[2]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((D*C))+~B*A*~((D*C))+~(~B)*A*(D*C)+~B*A*(D*C))"),
    .INIT(16'h5ccc))
    al_c35840ec (
    .a(al_9b9e072a),
    .b(al_ad4756a7[2]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1bc63bd7[2]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((D*~C))+~B*A*~((D*~C))+~(~B)*A*(D*~C)+~B*A*(D*~C))"),
    .INIT(16'hc5cc))
    al_b5961f1 (
    .a(al_9b9e072a),
    .b(al_ce7d4278[2]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_abc55d75[2]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((~D*~C))+~B*A*~((~D*~C))+~(~B)*A*(~D*~C)+~B*A*(~D*~C))"),
    .INIT(16'hccc5))
    al_4ccb051b (
    .a(al_9b9e072a),
    .b(al_47a64ed5[2]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_f8f25e7b[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_9f0224b3 (
    .a(al_1f23ce73[2]),
    .b(al_1bc63bd7[2]),
    .c(al_abc55d75[2]),
    .d(al_f8f25e7b[2]),
    .e(al_99c445b5[0]),
    .f(al_99c445b5[1]),
    .o(al_b6b411a2[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_d626c12a (
    .a(al_47a64ed5[3]),
    .b(al_75c1ef4c[3]),
    .c(al_ce7d4278[3]),
    .d(al_ad4756a7[3]),
    .e(al_879aba03[0]),
    .f(al_879aba03[1]),
    .o(al_a6b3d6e8));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)*~(A)+~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B*~(A)+~(~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*B*A+~(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B*A)"),
    .INIT(64'h7777722727722222))
    al_a625975b (
    .a(al_15b16fc6),
    .b(al_a6b3d6e8),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[3]),
    .f(al_75c0d27f[3]),
    .o(al_3ee9f2ae[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_b4faf18e (
    .a(al_3ee9f2ae[3]),
    .b(al_75c1ef4c[3]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1f23ce73[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_881766d2 (
    .a(al_3ee9f2ae[3]),
    .b(al_ad4756a7[3]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1bc63bd7[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_f5449418 (
    .a(al_3ee9f2ae[3]),
    .b(al_ce7d4278[3]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_abc55d75[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_8f9004c9 (
    .a(al_3ee9f2ae[3]),
    .b(al_47a64ed5[3]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_f8f25e7b[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_e15068f2 (
    .a(al_1f23ce73[3]),
    .b(al_1bc63bd7[3]),
    .c(al_abc55d75[3]),
    .d(al_f8f25e7b[3]),
    .e(al_99c445b5[0]),
    .f(al_99c445b5[1]),
    .o(al_b6b411a2[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_eae4d21b (
    .a(al_47a64ed5[4]),
    .b(al_75c1ef4c[4]),
    .c(al_ce7d4278[4]),
    .d(al_ad4756a7[4]),
    .e(al_879aba03[0]),
    .f(al_879aba03[1]),
    .o(al_518dbdc));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*(D@C))*~(B)*~(A)+~(E*(D@C))*B*~(A)+~(~(E*(D@C)))*B*A+~(E*(D@C))*B*A)"),
    .INIT(32'h27722222))
    al_5e0246f7 (
    .a(al_15b16fc6),
    .b(al_518dbdc),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[4]),
    .o(al_3ee9f2ae[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_e54efccf (
    .a(al_3ee9f2ae[4]),
    .b(al_75c1ef4c[4]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1f23ce73[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_3aef7788 (
    .a(al_3ee9f2ae[4]),
    .b(al_ad4756a7[4]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_1bc63bd7[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_a908c114 (
    .a(al_3ee9f2ae[4]),
    .b(al_ce7d4278[4]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_abc55d75[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_a31e6e4d (
    .a(al_3ee9f2ae[4]),
    .b(al_47a64ed5[4]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_f8f25e7b[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_e20905c8 (
    .a(al_1f23ce73[4]),
    .b(al_1bc63bd7[4]),
    .c(al_abc55d75[4]),
    .d(al_f8f25e7b[4]),
    .e(al_99c445b5[0]),
    .f(al_99c445b5[1]),
    .o(al_b6b411a2[4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_ef7a9585 (
    .a(al_7a00688b),
    .b(al_59addda8),
    .c(al_ac74f6f1),
    .d(al_80083fda[0]),
    .e(al_80083fda[1]),
    .o(al_a96c64c1));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    al_272ff7d6 (
    .a(al_891340a1),
    .b(al_a67dc86a[0]),
    .c(al_a67dc86a[1]),
    .d(al_c360bf4c[0]),
    .o(al_3f632af4));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h2c2f))
    al_a42eee81 (
    .a(al_891340a1),
    .b(al_a67dc86a[0]),
    .c(al_a67dc86a[1]),
    .d(al_e620c305),
    .o(al_94133c8a));
  AL_MAP_LUT6 #(
    .EQN("~((~D*~(~C*~(B*~A)))*~(E)*~(F)+(~D*~(~C*~(B*~A)))*E*~(F)+~((~D*~(~C*~(B*~A))))*E*F+(~D*~(~C*~(B*~A)))*E*F)"),
    .INIT(64'h0000ffffff0bff0b))
    al_56244be3 (
    .a(al_f0abb8e8[0]),
    .b(al_b4f15053),
    .c(al_fbbc76d0),
    .d(al_3f632af4),
    .e(al_94133c8a),
    .f(al_a67dc86a[2]),
    .o(al_c4e56ecb[0]));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~(~D*~(C*~(F*~(~B*~A)))))"),
    .INIT(64'hffff00efffff000f))
    al_d382b005 (
    .a(al_58fb4752[3]),
    .b(al_58fb4752[4]),
    .c(al_f7a41bbb),
    .d(al_a67dc86a[0]),
    .e(al_a67dc86a[1]),
    .f(al_df80405c),
    .o(al_fbbc76d0));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~(~D*~C*B*A))"),
    .INIT(64'hfff7000000000000))
    al_4eaaba07 (
    .a(al_99c9c113),
    .b(al_7a00688b),
    .c(al_80083fda[0]),
    .d(al_80083fda[1]),
    .e(al_6896ad14),
    .f(al_df80405c),
    .o(al_89c00c3));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(B*~(F*E*D*C)))"),
    .INIT(64'h5111111111111111))
    al_82c30d67 (
    .a(al_89c00c3),
    .b(al_a96c64c1),
    .c(al_93d3d349),
    .d(al_b5b02afa),
    .e(al_e71d5665),
    .f(al_e54eae62),
    .o(al_f0abb8e8[0]));
  AL_MAP_LUT6 #(
    .EQN("(F*~(E*D*C*B*A))"),
    .INIT(64'h7fffffff00000000))
    al_10c51201 (
    .a(al_93d3d349),
    .b(al_b5b02afa),
    .c(al_e71d5665),
    .d(al_e54eae62),
    .e(al_b6d031c2),
    .f(al_a67dc86a[0]),
    .o(al_b4f15053));
  AL_MAP_LUT6 #(
    .EQN("(F*A*~(E*D*C*B))"),
    .INIT(64'h2aaaaaaa00000000))
    al_261b112e (
    .a(al_a96c64c1),
    .b(al_93d3d349),
    .c(al_b5b02afa),
    .d(al_e71d5665),
    .e(al_e54eae62),
    .f(al_718bc19f),
    .o(al_28a9f919));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~A))*~(B)+D*(C*~A)*~(B)+~(D)*(C*~A)*B+D*(C*~A)*B)"),
    .INIT(16'h7340))
    al_d0137a55 (
    .a(al_891340a1),
    .b(al_a67dc86a[0]),
    .c(al_c360bf4c[0]),
    .d(al_90a0fe97[0]),
    .o(al_d03801fb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h03f0aaff03ffaaff))
    al_afcdfab9 (
    .a(al_d03801fb),
    .b(al_891340a1),
    .c(al_a67dc86a[0]),
    .d(al_a67dc86a[1]),
    .e(al_a67dc86a[2]),
    .f(al_e620c305),
    .o(al_634baaae));
  AL_MAP_LUT4 #(
    .EQN("~(C*~A*~(D*B))"),
    .INIT(16'hefaf))
    al_7f2e0fcd (
    .a(al_28a9f919),
    .b(al_aafc78b6),
    .c(al_634baaae),
    .d(al_718bc19f),
    .o(al_c4e56ecb[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F)"),
    .INIT(64'h13cf10cf13ff10ff))
    al_607ad5cd (
    .a(al_891340a1),
    .b(al_a67dc86a[0]),
    .c(al_a67dc86a[1]),
    .d(al_a67dc86a[2]),
    .e(al_e620c305),
    .f(al_90a0fe97[0]),
    .o(al_2873e816));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D*C*B))"),
    .INIT(16'hd555))
    al_e601e429 (
    .a(al_2873e816),
    .b(al_993745c8),
    .c(al_891340a1),
    .d(al_c360bf4c[0]),
    .o(al_c4e56ecb[2]));
  AL_MAP_LUT5 #(
    .EQN("((~B*A)*~(C)*~(D)*~(E)+(~B*A)*C*~(D)*~(E)+~((~B*A))*~(C)*D*~(E)+(~B*A)*~(C)*D*~(E)+~((~B*A))*C*~(D)*E+(~B*A)*C*~(D)*E+~((~B*A))*~(C)*D*E+(~B*A)*~(C)*D*E+~((~B*A))*C*D*E+(~B*A)*C*D*E)"),
    .INIT(32'hfff00f22))
    al_23b1c603 (
    .a(al_74e913f6),
    .b(al_2bb5f88f),
    .c(al_1e3dbb5f),
    .d(al_c46598af[0]),
    .e(al_c46598af[1]),
    .o(al_7c5b4e5e[0]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(~C*B*A))"),
    .INIT(16'hff08))
    al_992cfeac (
    .a(al_74e913f6),
    .b(al_2bb5f88f),
    .c(al_c46598af[0]),
    .d(al_c46598af[1]),
    .o(al_7c5b4e5e[1]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_c72a60d2 (
    .a(al_97784c51),
    .b(al_1e500c02),
    .c(al_25aa754),
    .o(al_98c339b0));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_14048e58 (
    .a(al_9fcbbf12),
    .b(al_1e500c02),
    .c(al_25aa754),
    .o(al_8ee904a8));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_6780f75a (
    .a(al_a4d81981),
    .b(al_1e500c02),
    .c(al_25aa754),
    .o(al_62952198));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_313e0559 (
    .a(al_cf11b78b[0]),
    .b(al_a67dc86a[0]),
    .c(al_a67dc86a[1]),
    .d(al_a67dc86a[2]),
    .e(al_898823b1),
    .o(al_1e500c02));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_64d6f15d (
    .a(al_d3154fbb),
    .b(al_1e500c02),
    .c(al_25aa754),
    .o(al_92e98f85));
  AL_DFF_0 al_e66edca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_456c110a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_58ef9f1a));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_fd5d0b41 (
    .a(al_ebce8257),
    .b(al_456c110a),
    .o(al_81e393a7));
  AL_DFF_0 al_62ecacfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_81e393a7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45b542b0));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_ebf242c1 (
    .a(al_45b542b0),
    .b(al_456c110a),
    .o(al_b79e57b1));
  AL_DFF_0 al_29ae1406 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b79e57b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fa36ca4c));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_7199e529 (
    .a(al_fa36ca4c),
    .b(al_456c110a),
    .o(al_1358b03f));
  AL_DFF_0 al_90de0a0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1358b03f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49c007fc));
  AL_DFF_0 al_83d85781 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_648bb7aa),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_ebce8257));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    al_15d81b01 (
    .a(al_ebce8257),
    .b(al_456c110a),
    .c(al_4b38e0f3),
    .o(al_648bb7aa));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_fb6bb359 (
    .a(al_648bb7aa),
    .b(al_ebce8257),
    .c(al_898823b1),
    .o(al_afe8fb08));
  AL_DFF_0 al_fcf056d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_afe8fb08),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2d3f245b));
  AL_DFF_0 al_571bb883 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff3a70dc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c104e46));
  AL_DFF_0 al_655c7db4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d76e6af),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_c56a3e50));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    al_27d07ea1 (
    .a(al_28a9f919),
    .b(al_c56a3e50),
    .c(al_90a0fe97[0]),
    .o(al_4d76e6af));
  AL_DFF_0 al_449f2a40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5d5ab475[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_cfaa4b74));
  AL_DFF_0 al_a90503db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5d5ab475[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_1c7e0f23));
  AL_DFF_0 al_e2108b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5d5ab475[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_80cba1f));
  AL_DFF_0 al_108202ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5d5ab475[3]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2f87218f));
  AL_DFF_0 al_a90efe94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5d5ab475[4]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2d60bf7c));
  AL_DFF_0 al_d5aa1cbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b5844352[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_1fe24196));
  AL_DFF_0 al_aff5ebca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b5844352[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_4c2bab56));
  AL_DFF_0 al_ed50d62f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b5844352[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b325b551));
  AL_DFF_0 al_38f520af (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b5844352[3]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2761bf91));
  AL_DFF_0 al_d7f70db0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a65f5154[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_a5d3389d));
  AL_DFF_0 al_bf58e226 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a65f5154[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_840aa4cd));
  AL_DFF_0 al_4ac3e22b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a65f5154[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_6e2c4231));
  AL_DFF_0 al_d87bc111 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a65f5154[3]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_af3006e2));
  AL_DFF_0 al_2e955ed7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56b3021d[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_6cdb74d6));
  AL_DFF_0 al_98b5eedc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56b3021d[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_6ab92c75));
  AL_DFF_0 al_a147ea40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56b3021d[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_287c07f8));
  AL_DFF_0 al_6dddf73f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56b3021d[3]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_f9b2e036));
  AL_DFF_0 al_a6861000 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf91271d[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_5341a91c));
  AL_DFF_0 al_65447aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf91271d[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_591ab1d4));
  AL_DFF_0 al_65b5ddb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf91271d[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b23d9425));
  AL_DFF_0 al_90cc7a2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf91271d[3]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_a02f02e8));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_bf859581 (
    .a(al_a67dc86a[0]),
    .b(al_a67dc86a[1]),
    .c(al_a67dc86a[2]),
    .o(al_993745c8));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_54ce817 (
    .a(al_993745c8),
    .b(al_b93da8d5[0]),
    .c(al_b93da8d5[1]),
    .o(al_9fcbbf12));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5d40aeca (
    .a(al_9fcbbf12),
    .b(al_c360bf4c[0]),
    .o(al_c00d3bb));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_72350952 (
    .a(al_c00d3bb),
    .b(al_a5d3389d),
    .c(al_840aa4cd),
    .d(al_6e2c4231),
    .e(al_af3006e2),
    .f(al_d2824414),
    .o(al_a65f5154[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_49dc4959 (
    .a(al_c00d3bb),
    .b(al_a5d3389d),
    .c(al_d2824414),
    .o(al_a65f5154[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_39f46385 (
    .a(al_c00d3bb),
    .b(al_a5d3389d),
    .c(al_840aa4cd),
    .d(al_d2824414),
    .o(al_a65f5154[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_a23b47c0 (
    .a(al_c00d3bb),
    .b(al_a5d3389d),
    .c(al_840aa4cd),
    .d(al_6e2c4231),
    .e(al_d2824414),
    .o(al_a65f5154[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_458e4cff (
    .a(al_993745c8),
    .b(al_b93da8d5[0]),
    .c(al_b93da8d5[1]),
    .o(al_a4d81981));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_7c2efa94 (
    .a(al_a4d81981),
    .b(al_c360bf4c[0]),
    .o(al_69a88833));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_80e74ad9 (
    .a(al_69a88833),
    .b(al_6cdb74d6),
    .c(al_6ab92c75),
    .d(al_287c07f8),
    .e(al_f9b2e036),
    .f(al_7cad9721),
    .o(al_56b3021d[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_476c9844 (
    .a(al_69a88833),
    .b(al_6cdb74d6),
    .c(al_7cad9721),
    .o(al_56b3021d[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_5367b864 (
    .a(al_69a88833),
    .b(al_6cdb74d6),
    .c(al_6ab92c75),
    .d(al_7cad9721),
    .o(al_56b3021d[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_6fb8d36b (
    .a(al_69a88833),
    .b(al_6cdb74d6),
    .c(al_6ab92c75),
    .d(al_287c07f8),
    .e(al_7cad9721),
    .o(al_56b3021d[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_7f43bc5c (
    .a(al_993745c8),
    .b(al_b93da8d5[0]),
    .c(al_b93da8d5[1]),
    .o(al_d3154fbb));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_cb4144ba (
    .a(al_d3154fbb),
    .b(al_c360bf4c[0]),
    .o(al_9d7e8bc9));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_8bf31ca9 (
    .a(al_9d7e8bc9),
    .b(al_5341a91c),
    .c(al_591ab1d4),
    .d(al_b23d9425),
    .e(al_a02f02e8),
    .f(al_681e3ff2),
    .o(al_cf91271d[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_4aed98ea (
    .a(al_9d7e8bc9),
    .b(al_5341a91c),
    .c(al_681e3ff2),
    .o(al_cf91271d[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_74745181 (
    .a(al_9d7e8bc9),
    .b(al_5341a91c),
    .c(al_591ab1d4),
    .d(al_681e3ff2),
    .o(al_cf91271d[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_2a41fe7f (
    .a(al_9d7e8bc9),
    .b(al_5341a91c),
    .c(al_591ab1d4),
    .d(al_b23d9425),
    .e(al_681e3ff2),
    .o(al_cf91271d[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_de08dc00 (
    .a(al_993745c8),
    .b(al_b93da8d5[0]),
    .c(al_b93da8d5[1]),
    .o(al_97784c51));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_e0384135 (
    .a(al_97784c51),
    .b(al_c360bf4c[0]),
    .o(al_e7604954));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_65f5efee (
    .a(al_e7604954),
    .b(al_1fe24196),
    .c(al_4c2bab56),
    .d(al_b325b551),
    .e(al_2761bf91),
    .f(al_280c0ef0),
    .o(al_b5844352[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_fb16c109 (
    .a(al_e7604954),
    .b(al_1fe24196),
    .c(al_280c0ef0),
    .o(al_b5844352[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_6dd96c12 (
    .a(al_e7604954),
    .b(al_1fe24196),
    .c(al_4c2bab56),
    .d(al_280c0ef0),
    .o(al_b5844352[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_a78bb49d (
    .a(al_e7604954),
    .b(al_1fe24196),
    .c(al_4c2bab56),
    .d(al_b325b551),
    .e(al_280c0ef0),
    .o(al_b5844352[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_7e2048b (
    .a(al_a65f5154[3]),
    .b(al_a65f5154[0]),
    .c(al_a65f5154[1]),
    .d(al_a65f5154[2]),
    .o(al_c2faf058[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_48bc98e4 (
    .a(al_56b3021d[3]),
    .b(al_56b3021d[0]),
    .c(al_56b3021d[1]),
    .d(al_56b3021d[2]),
    .o(al_c2faf058[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_635a7d8a (
    .a(al_cf91271d[3]),
    .b(al_cf91271d[0]),
    .c(al_cf91271d[1]),
    .d(al_cf91271d[2]),
    .o(al_c2faf058[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_c562717e (
    .a(al_b5844352[3]),
    .b(al_b5844352[0]),
    .c(al_b5844352[1]),
    .d(al_b5844352[2]),
    .o(al_c2faf058[0]));
  AL_DFF_0 al_2e581ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c2faf058[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_280c0ef0));
  AL_DFF_0 al_495ffa0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c2faf058[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d2824414));
  AL_DFF_0 al_d7462e02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c2faf058[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cad9721));
  AL_DFF_0 al_39f68928 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c2faf058[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_681e3ff2));
  AL_DFF_0 al_2b32b67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f9833848),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18326672));
  AL_DFF_0 al_44546ccb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[24]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_688aeb95));
  AL_DFF_0 al_42e339ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[25]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_8cae5877));
  AL_DFF_0 al_d2e791c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[26]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_e769a1ac));
  AL_DFF_0 al_bfb16e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[27]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_a4dd8227));
  AL_DFF_0 al_c1cd9d61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[28]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_da2e6045));
  AL_DFF_0 al_1b8bfc22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[29]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_ac3b1637));
  AL_DFF_0 al_bfbfc5b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[30]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_533b1c82));
  AL_DFF_0 al_eba4faa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[31]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_41ef913c));
  AL_DFF_0 al_10f18eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[32]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_17bf017e));
  AL_DFF_0 al_76b6532b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[33]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_c952c11c));
  AL_DFF_0 al_a08fc634 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[34]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_ac45c87a));
  AL_DFF_0 al_d6c427d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[35]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_83d9c8d2));
  AL_DFF_0 al_7477445b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[36]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_227f8a62));
  AL_DFF_0 al_c237cdee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[37]),
    .en(al_98c339b0),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_4d37ff05));
  AL_DFF_0 al_1b0f1ace (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d38737b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5ec2c98e));
  AL_DFF_0 al_39af5fdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[24]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_bbfb7745));
  AL_DFF_0 al_96691900 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[25]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_f71dba21));
  AL_DFF_0 al_dd9de9d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[26]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_267ffb9b));
  AL_DFF_0 al_576b466f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[27]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_97814ee2));
  AL_DFF_0 al_7afd1148 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[28]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2b60c4d7));
  AL_DFF_0 al_d5a17f2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[29]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_f9500eb2));
  AL_DFF_0 al_1beeea65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[30]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_85770a25));
  AL_DFF_0 al_8ce041b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[31]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_457533f2));
  AL_DFF_0 al_311f4903 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[32]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_5f86f74e));
  AL_DFF_0 al_1019741e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[33]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_e5cd290d));
  AL_DFF_0 al_3aa107d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[34]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2f21552f));
  AL_DFF_0 al_c4702e1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[35]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_232e33c9));
  AL_DFF_0 al_95dc1e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[36]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_c8afcceb));
  AL_DFF_0 al_cae8563f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[37]),
    .en(al_8ee904a8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_50f5aee2));
  AL_DFF_0 al_f52b7df0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_640fb7ec),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_370aa1bb));
  AL_DFF_0 al_a3ae0a94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[24]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_1b8721f8));
  AL_DFF_0 al_c1686ad6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[25]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_1f70c9fe));
  AL_DFF_0 al_6d89dd64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[26]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9e92954d));
  AL_DFF_0 al_e4c7aee1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[27]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_736e37f2));
  AL_DFF_0 al_674a19fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[28]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_4f668848));
  AL_DFF_0 al_51ef5178 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[29]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9cb32c9b));
  AL_DFF_0 al_409d8357 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[30]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_899fc7f2));
  AL_DFF_0 al_fe1c45e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[31]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_e9f106ba));
  AL_DFF_0 al_91421113 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[32]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_fd00fe9e));
  AL_DFF_0 al_2d7ad1a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[33]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_1f4c68e6));
  AL_DFF_0 al_b39d80d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[34]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d17a0773));
  AL_DFF_0 al_1eb2e263 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[35]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_95538c25));
  AL_DFF_0 al_895955d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[36]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_e0aa83ea));
  AL_DFF_0 al_67e86cbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[37]),
    .en(al_62952198),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_c5c92715));
  AL_DFF_0 al_29e27edb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a315f23),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_72b4a28e));
  AL_DFF_0 al_168a559b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[24]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b741880));
  AL_DFF_0 al_8f941f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[25]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d177c6b8));
  AL_DFF_0 al_9136680d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[26]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_bf6feeb3));
  AL_DFF_0 al_cd541dd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[27]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_f31ca00d));
  AL_DFF_0 al_9c7737dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[28]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_37cdc8a1));
  AL_DFF_0 al_fddb7f40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[29]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_8ff2e306));
  AL_DFF_0 al_4196640b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[30]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_993b1b0f));
  AL_DFF_0 al_1b5b0b6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[31]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_bc420de3));
  AL_DFF_0 al_f4fb4927 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[32]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_ece57492));
  AL_DFF_0 al_4ad9c5b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[33]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_3c73e97d));
  AL_DFF_0 al_145559c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[34]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_3b11a186));
  AL_DFF_0 al_d0eda2c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[35]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b0e11bf3));
  AL_DFF_0 al_5653bcc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[36]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9f6af9ba));
  AL_DFF_0 al_92613911 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[37]),
    .en(al_92e98f85),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_c7421999));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_c6df0239 (
    .a(al_9fcbbf12),
    .b(al_1e500c02),
    .c(al_5ec2c98e),
    .d(al_25aa754),
    .e(al_3ee0d55a),
    .o(al_4d38737b));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_76950a8a (
    .a(al_97784c51),
    .b(al_1e500c02),
    .c(al_18326672),
    .d(al_25aa754),
    .e(al_3ee0d55a),
    .o(al_f9833848));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_6f467658 (
    .a(al_d3154fbb),
    .b(al_1e500c02),
    .c(al_72b4a28e),
    .d(al_25aa754),
    .e(al_3ee0d55a),
    .o(al_a315f23));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_42eabf7e (
    .a(al_a4d81981),
    .b(al_1e500c02),
    .c(al_370aa1bb),
    .d(al_25aa754),
    .e(al_3ee0d55a),
    .o(al_640fb7ec));
  AL_DFF_0 al_c860efcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d549f91e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25aa754));
  AL_DFF_0 al_c29214b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d7619b2[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2b3c55e4));
  AL_DFF_0 al_f5d9a287 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c84bba78),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_1c1fb07a));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_956ab1ac (
    .a(al_da34749d),
    .b(al_71f78ff1[46]),
    .c(al_c46598af[0]),
    .d(al_c46598af[1]),
    .o(al_d102b3df));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~(B*A)))"),
    .INIT(16'h0f08))
    al_83cdb984 (
    .a(al_74e913f6),
    .b(al_d102b3df),
    .c(al_1e3dbb5f),
    .d(al_1c1fb07a),
    .o(al_c84bba78));
  AL_DFF_0 al_59a983cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d42c904d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf11b78b[0]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_d2d2a291 (
    .a(al_8a415a42),
    .b(al_6896ad14),
    .c(al_a67dc86a[0]),
    .d(al_a67dc86a[1]),
    .e(al_a67dc86a[2]),
    .o(al_d42c904d));
  AL_DFF_0 al_921ecbe5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_898823b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c9229ee));
  AL_DFF_0 al_c81abdc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c9229ee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6e223da));
  AL_DFF_0 al_fab36d83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6e223da),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e1f18395));
  AL_DFF_0 al_8c6372c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1f18395),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6896ad14));
  AL_DFF_0 al_f5bfc17c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_53b2015),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbeafa67[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    al_4f1b2398 (
    .a(al_28a9f919),
    .b(al_cbeafa67[0]),
    .c(al_b93da8d5[2]),
    .d(al_3ee0d55a),
    .o(al_53b2015));
  AL_DFF_0 al_59c6f360 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_31adf876[0]));
  AL_DFF_0 al_626152f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_31adf876[1]));
  AL_DFF_0 al_e135206b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d76fa964[0]));
  AL_DFF_0 al_e7f2fdf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c4e56ecb[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_a67dc86a[0]));
  AL_DFF_0 al_be3c0f1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c4e56ecb[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_a67dc86a[1]));
  AL_DFF_0 al_84e2ac82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c4e56ecb[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_a67dc86a[2]));
  AL_DFF_0 al_46864a06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c5b4e5e[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_c46598af[0]));
  AL_DFF_0 al_d0d3e20b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c5b4e5e[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_c46598af[1]));
  AL_DFF_0 al_128dc602 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[0]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[0]));
  AL_DFF_0 al_efa394e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[1]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[1]));
  AL_DFF_0 al_2b47b63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[2]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[2]));
  AL_DFF_0 al_a12a64dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[11]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[11]));
  AL_DFF_0 al_10708ebe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[12]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[12]));
  AL_DFF_0 al_d50b5838 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[13]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[13]));
  AL_DFF_0 al_673117df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[14]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[14]));
  AL_DFF_0 al_c7bb80a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[15]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[15]));
  AL_DFF_0 al_5f048f58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[16]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[16]));
  AL_DFF_0 al_5f47eca5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[17]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[17]));
  AL_DFF_0 al_8726eaf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[24]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[24]));
  AL_DFF_0 al_9c9606a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[25]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[25]));
  AL_DFF_0 al_8b1b433e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[26]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[26]));
  AL_DFF_0 al_987ca071 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[27]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[27]));
  AL_DFF_0 al_e3c6f598 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[28]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[28]));
  AL_DFF_0 al_fca371bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[29]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[29]));
  AL_DFF_0 al_34dbbcce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[30]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[30]));
  AL_DFF_0 al_2fd2dac1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[31]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[31]));
  AL_DFF_0 al_50dfafcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[32]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[32]));
  AL_DFF_0 al_8d98e004 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[33]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[33]));
  AL_DFF_0 al_c5d37243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[34]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[34]));
  AL_DFF_0 al_90a7cdbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[35]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[35]));
  AL_DFF_0 al_d6af8aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[36]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[36]));
  AL_DFF_0 al_6b602d75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[37]),
    .en(al_52665bb8),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_58851aab[37]));
  AL_DFF_0 al_e3a12c74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f8f25e7b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_47a64ed5[0]));
  AL_DFF_0 al_b9f1d768 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f8f25e7b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_47a64ed5[1]));
  AL_DFF_0 al_c304891 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f8f25e7b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_47a64ed5[2]));
  AL_DFF_0 al_d1645bdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f8f25e7b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_47a64ed5[3]));
  AL_DFF_0 al_138fe171 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f8f25e7b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_47a64ed5[4]));
  AL_DFF_0 al_a5b6c6fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f23ce73[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75c1ef4c[0]));
  AL_DFF_0 al_4ab97fb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f23ce73[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75c1ef4c[1]));
  AL_DFF_0 al_9e30742e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f23ce73[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75c1ef4c[2]));
  AL_DFF_0 al_d2517ba5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f23ce73[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75c1ef4c[3]));
  AL_DFF_0 al_dbc1dffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f23ce73[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75c1ef4c[4]));
  AL_DFF_0 al_1ffc754 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_abc55d75[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce7d4278[0]));
  AL_DFF_0 al_690a6aa2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_abc55d75[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce7d4278[1]));
  AL_DFF_0 al_e595e886 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_abc55d75[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce7d4278[2]));
  AL_DFF_0 al_79e6bc3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_abc55d75[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce7d4278[3]));
  AL_DFF_0 al_dc633b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_abc55d75[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce7d4278[4]));
  AL_DFF_0 al_7c1c4ca9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1bc63bd7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad4756a7[0]));
  AL_DFF_0 al_f217dd79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1bc63bd7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad4756a7[1]));
  AL_DFF_0 al_dc3aa3df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1bc63bd7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad4756a7[2]));
  AL_DFF_0 al_6521d010 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1bc63bd7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad4756a7[3]));
  AL_DFF_0 al_59d48528 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1bc63bd7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad4756a7[4]));
  AL_DFF_0 al_27c50c69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7711fc3[3]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_81f91ff1[3]));
  AL_DFF_0 al_c51f1efa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7711fc3[4]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_81f91ff1[4]));
  AL_DFF_0 al_de8b4ad4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7711fc3[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_81f91ff1[0]));
  AL_DFF_0 al_b2584495 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7711fc3[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_81f91ff1[1]));
  AL_DFF_0 al_5ec6f5df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7711fc3[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_81f91ff1[2]));
  AL_DFF_0 al_630b625 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[0]));
  AL_DFF_0 al_457da81c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[1]));
  AL_DFF_0 al_d74f27fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[2]));
  AL_DFF_0 al_6ce3dde4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[11]));
  AL_DFF_0 al_56d5ba37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[12]));
  AL_DFF_0 al_5cd52c94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[13]));
  AL_DFF_0 al_6ce1da39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[14]));
  AL_DFF_0 al_900a24bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[15]));
  AL_DFF_0 al_8271e6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[16]));
  AL_DFF_0 al_85d35ca2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[17]));
  AL_DFF_0 al_8a966314 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[24]));
  AL_DFF_0 al_416b73bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[25]));
  AL_DFF_0 al_26b11d63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[26]));
  AL_DFF_0 al_2b2804bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[27]));
  AL_DFF_0 al_ac62aa32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[28]));
  AL_DFF_0 al_fe57193e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[29]));
  AL_DFF_0 al_12c93e7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[30]));
  AL_DFF_0 al_3b9358f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[31]));
  AL_DFF_0 al_c28e2b62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[32]));
  AL_DFF_0 al_f443b518 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[33]));
  AL_DFF_0 al_7c366d06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[34]));
  AL_DFF_0 al_53b29fcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[35]));
  AL_DFF_0 al_aca53f2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[36]));
  AL_DFF_0 al_face12e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[37]));
  AL_DFF_0 al_f3e08773 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[44]));
  AL_DFF_0 al_8a8ef2f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[45]));
  AL_DFF_0 al_add45e14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[46]));
  AL_DFF_0 al_3c03efba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6be20a95[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b93da8d5[48]));
  AL_DFF_0 al_45f76bad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[0]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[0]));
  AL_DFF_0 al_c8d97ecb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[1]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[1]));
  AL_DFF_0 al_50550b2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[2]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[2]));
  AL_DFF_0 al_27f58777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[11]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[11]));
  AL_DFF_0 al_29c86684 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[12]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[12]));
  AL_DFF_0 al_bd8b8139 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[13]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[13]));
  AL_DFF_0 al_96d79109 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[14]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[14]));
  AL_DFF_0 al_212349fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[15]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[15]));
  AL_DFF_0 al_ef389046 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[16]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[16]));
  AL_DFF_0 al_83996c7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[17]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[17]));
  AL_DFF_0 al_7be85095 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[24]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[24]));
  AL_DFF_0 al_2cfccfa5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[25]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[25]));
  AL_DFF_0 al_68e7cc91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[26]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[26]));
  AL_DFF_0 al_3409fc64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[27]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[27]));
  AL_DFF_0 al_b69be5da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[28]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[28]));
  AL_DFF_0 al_83670acb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[29]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[29]));
  AL_DFF_0 al_cc1c9845 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[30]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[30]));
  AL_DFF_0 al_776d994d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[31]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[31]));
  AL_DFF_0 al_dd5e22b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[32]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[32]));
  AL_DFF_0 al_cd282574 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[33]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[33]));
  AL_DFF_0 al_556251da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[34]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[34]));
  AL_DFF_0 al_96abff62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[35]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[35]));
  AL_DFF_0 al_6efdaae1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[36]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[36]));
  AL_DFF_0 al_94f01071 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[37]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[37]));
  AL_DFF_0 al_b788adb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[44]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[44]));
  AL_DFF_0 al_547a07d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[45]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[45]));
  AL_DFF_0 al_c865ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[46]),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[46]));
  AL_DFF_0 al_d513d097 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4ecf439),
    .en(al_5453b759[0]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_77634075[48]));
  AL_DFF_0 al_72c27c4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[0]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[0]));
  AL_DFF_0 al_c67210a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[1]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[1]));
  AL_DFF_0 al_26fb132d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[2]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[2]));
  AL_DFF_0 al_94945c79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[11]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[11]));
  AL_DFF_0 al_93ce133c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[12]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[12]));
  AL_DFF_0 al_6308ef0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[13]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[13]));
  AL_DFF_0 al_1bf005 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[14]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[14]));
  AL_DFF_0 al_6f9a5b9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[15]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[15]));
  AL_DFF_0 al_47242d8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[16]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[16]));
  AL_DFF_0 al_89cc2ba0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[17]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[17]));
  AL_DFF_0 al_a66c1388 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[24]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[24]));
  AL_DFF_0 al_4fc56c41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[25]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[25]));
  AL_DFF_0 al_8415064a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[26]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[26]));
  AL_DFF_0 al_2d6cf803 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[27]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[27]));
  AL_DFF_0 al_3f151a57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[28]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[28]));
  AL_DFF_0 al_64f3e113 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[29]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[29]));
  AL_DFF_0 al_bc1ede32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[30]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[30]));
  AL_DFF_0 al_f2bb15f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[31]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[31]));
  AL_DFF_0 al_28cd1607 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[32]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[32]));
  AL_DFF_0 al_ac11ca34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[33]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[33]));
  AL_DFF_0 al_5bb0e84d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[34]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[34]));
  AL_DFF_0 al_55f07844 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[35]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[35]));
  AL_DFF_0 al_e16bdae9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[36]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[36]));
  AL_DFF_0 al_e8af5de8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[37]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[37]));
  AL_DFF_0 al_1f73557f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[44]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[44]));
  AL_DFF_0 al_6eadd7eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[45]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[45]));
  AL_DFF_0 al_283c9b50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[46]),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[46]));
  AL_DFF_0 al_b0684a93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4ecf439),
    .en(al_5453b759[1]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_b9ba8b6c[48]));
  AL_DFF_0 al_4f2808e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[0]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[0]));
  AL_DFF_0 al_4c6d390a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[1]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[1]));
  AL_DFF_0 al_1980d79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[2]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[2]));
  AL_DFF_0 al_673c6318 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[11]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[11]));
  AL_DFF_0 al_c202155e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[12]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[12]));
  AL_DFF_0 al_d5b23716 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[13]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[13]));
  AL_DFF_0 al_a5bfd85d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[14]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[14]));
  AL_DFF_0 al_772a326d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[15]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[15]));
  AL_DFF_0 al_d81ae086 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[16]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[16]));
  AL_DFF_0 al_12ce4854 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[17]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[17]));
  AL_DFF_0 al_ce4330c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[24]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[24]));
  AL_DFF_0 al_60203319 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[25]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[25]));
  AL_DFF_0 al_96bd10a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[26]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[26]));
  AL_DFF_0 al_1b80b1e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[27]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[27]));
  AL_DFF_0 al_be8b6bf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[28]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[28]));
  AL_DFF_0 al_d96a812e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[29]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[29]));
  AL_DFF_0 al_2b1205bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[30]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[30]));
  AL_DFF_0 al_b7a7cf5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[31]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[31]));
  AL_DFF_0 al_43c1e8a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[32]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[32]));
  AL_DFF_0 al_c521b1e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[33]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[33]));
  AL_DFF_0 al_9de2317d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[34]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[34]));
  AL_DFF_0 al_aa54279 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[35]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[35]));
  AL_DFF_0 al_f1a53502 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[36]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[36]));
  AL_DFF_0 al_2354346b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[37]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[37]));
  AL_DFF_0 al_b0b3543f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[44]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[44]));
  AL_DFF_0 al_5ee7bc1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[45]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[45]));
  AL_DFF_0 al_42d7710a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[46]),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[46]));
  AL_DFF_0 al_378da6a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4ecf439),
    .en(al_5453b759[2]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_9c434c4a[48]));
  AL_DFF_0 al_bb27b51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[0]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[0]));
  AL_DFF_0 al_5aecbe95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[1]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[1]));
  AL_DFF_0 al_44dfdc7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[2]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[2]));
  AL_DFF_0 al_cbf33a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[11]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[11]));
  AL_DFF_0 al_a489be44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[12]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[12]));
  AL_DFF_0 al_4c965540 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[13]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[13]));
  AL_DFF_0 al_dd9b0b50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[14]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[14]));
  AL_DFF_0 al_78a47434 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[15]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[15]));
  AL_DFF_0 al_898219ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[16]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[16]));
  AL_DFF_0 al_d3209906 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[17]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[17]));
  AL_DFF_0 al_ce217a1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[24]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[24]));
  AL_DFF_0 al_c4e2cf12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[25]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[25]));
  AL_DFF_0 al_733a0b99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[26]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[26]));
  AL_DFF_0 al_b0bd031c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[27]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[27]));
  AL_DFF_0 al_a66e39a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[28]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[28]));
  AL_DFF_0 al_610b2be3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[29]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[29]));
  AL_DFF_0 al_f36abe5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[30]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[30]));
  AL_DFF_0 al_b8577da8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[31]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[31]));
  AL_DFF_0 al_8227babf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[32]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[32]));
  AL_DFF_0 al_284802ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[33]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[33]));
  AL_DFF_0 al_9ddc3138 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[34]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[34]));
  AL_DFF_0 al_413b723d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[35]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[35]));
  AL_DFF_0 al_ba86f6dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[36]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[36]));
  AL_DFF_0 al_7884aad2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[37]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[37]));
  AL_DFF_0 al_c4f86691 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[44]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[44]));
  AL_DFF_0 al_a101ef2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[45]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[45]));
  AL_DFF_0 al_9b5bd507 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e489598[46]),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[46]));
  AL_DFF_0 al_6d0a8b2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4ecf439),
    .en(al_5453b759[3]),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_d3350acc[48]));
  AL_DFF_0 al_f21ef0ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_765e8240[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_99c445b5[0]));
  AL_DFF_0 al_601d2be6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_765e8240[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_99c445b5[1]));
  AL_DFF_0 al_f2bedc8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e484293d[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_879aba03[0]));
  AL_DFF_0 al_43b25347 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e484293d[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_879aba03[1]));
  AL_DFF_0 al_a22ac0fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[0]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2a06982[0]));
  AL_DFF_0 al_54a26985 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[1]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2a06982[1]));
  AL_DFF_0 al_fd7fe027 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[2]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2a06982[2]));
  AL_DFF_0 al_b1d7a8b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[3]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2a06982[3]));
  AL_DFF_0 al_4a1a8977 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[4]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2a06982[4]));
  AL_DFF_0 al_49289ed7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[0]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c3bcd0f7[0]));
  AL_DFF_0 al_9ab1eb99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[1]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c3bcd0f7[1]));
  AL_DFF_0 al_cc4d39f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[2]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c3bcd0f7[2]));
  AL_DFF_0 al_abe5f793 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[3]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c3bcd0f7[3]));
  AL_DFF_0 al_b58ccdbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[4]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c3bcd0f7[4]));
  AL_DFF_0 al_78b1e4a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[0]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35348eec[0]));
  AL_DFF_0 al_4cb62166 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[1]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35348eec[1]));
  AL_DFF_0 al_6c91276e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[2]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35348eec[2]));
  AL_DFF_0 al_cce70084 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[3]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35348eec[3]));
  AL_DFF_0 al_caa51c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[4]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35348eec[4]));
  AL_DFF_0 al_52533aef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[0]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd4b89ad[0]));
  AL_DFF_0 al_e87ae80d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[1]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd4b89ad[1]));
  AL_DFF_0 al_39ea17c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[2]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd4b89ad[2]));
  AL_DFF_0 al_11b6498c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[3]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd4b89ad[3]));
  AL_DFF_0 al_42610eb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6b411a2[4]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd4b89ad[4]));
  AL_DFF_0 al_e93e2526 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d5c3e265[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_ffbe21a4[0]));
  AL_DFF_0 al_8cdeb9c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d5c3e265[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_ffbe21a4[1]));
  AL_DFF_0 al_d90a5a3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_845e0bd1[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_73f8a8a7[0]));
  AL_DFF_0 al_3c585793 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_845e0bd1[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_73f8a8a7[1]));
  AL_DFF_0 al_edb06633 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_845e0bd1[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_73f8a8a7[2]));
  AL_DFF_0 al_bc7440af (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_845e0bd1[3]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_73f8a8a7[3]));
  AL_DFF_0 al_3b8bc595 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[0]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[0]));
  AL_DFF_0 al_c4be6dce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[1]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[1]));
  AL_DFF_0 al_90aacb0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[2]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[2]));
  AL_DFF_0 al_c1210943 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[11]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[11]));
  AL_DFF_0 al_c3573a39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[12]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[12]));
  AL_DFF_0 al_59b0a7b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[13]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[13]));
  AL_DFF_0 al_d4e54599 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[14]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[14]));
  AL_DFF_0 al_9abba269 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[15]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[15]));
  AL_DFF_0 al_90495b7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[16]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[16]));
  AL_DFF_0 al_ea33f5cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[17]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[17]));
  AL_DFF_0 al_da7fa244 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[44]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[44]));
  AL_DFF_0 al_a78eeff8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[45]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[45]));
  AL_DFF_0 al_7da4321d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[46]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[46]));
  AL_DFF_0 al_69426746 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[48]),
    .en(al_10206333[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0482f12[48]));
  AL_DFF_0 al_b9c55779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[0]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[0]));
  AL_DFF_0 al_99b48953 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[1]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[1]));
  AL_DFF_0 al_b3eb530 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[2]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[2]));
  AL_DFF_0 al_67aebb35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[11]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[11]));
  AL_DFF_0 al_3c25454d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[12]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[12]));
  AL_DFF_0 al_bf3a40fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[13]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[13]));
  AL_DFF_0 al_9178e299 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[14]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[14]));
  AL_DFF_0 al_9fa9e892 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[15]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[15]));
  AL_DFF_0 al_4b0e86b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[16]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[16]));
  AL_DFF_0 al_6864254e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[17]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[17]));
  AL_DFF_0 al_22efe9b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[44]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[44]));
  AL_DFF_0 al_1ade5382 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[45]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[45]));
  AL_DFF_0 al_5325022b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[46]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[46]));
  AL_DFF_0 al_33af9aee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[48]),
    .en(al_10206333[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b620bb0[48]));
  AL_DFF_0 al_3dcae609 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[0]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[0]));
  AL_DFF_0 al_6aa31eaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[1]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[1]));
  AL_DFF_0 al_dc6f3152 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[2]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[2]));
  AL_DFF_0 al_14167067 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[11]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[11]));
  AL_DFF_0 al_ea548761 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[12]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[12]));
  AL_DFF_0 al_50132da0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[13]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[13]));
  AL_DFF_0 al_2c658733 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[14]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[14]));
  AL_DFF_0 al_6f7788c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[15]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[15]));
  AL_DFF_0 al_f416ca2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[16]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[16]));
  AL_DFF_0 al_e4ac636f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[17]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[17]));
  AL_DFF_0 al_d754f989 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[44]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[44]));
  AL_DFF_0 al_46c0f460 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[45]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[45]));
  AL_DFF_0 al_37188614 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[46]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[46]));
  AL_DFF_0 al_f0ce4fd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[48]),
    .en(al_10206333[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5104c4f[48]));
  AL_DFF_0 al_68ef07b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[0]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[0]));
  AL_DFF_0 al_4efa59bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[1]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[1]));
  AL_DFF_0 al_b9591cba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[2]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[2]));
  AL_DFF_0 al_943226c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[11]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[11]));
  AL_DFF_0 al_4a95b10d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[12]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[12]));
  AL_DFF_0 al_7395efa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[13]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[13]));
  AL_DFF_0 al_5527974d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[14]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[14]));
  AL_DFF_0 al_3e629cda (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[15]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[15]));
  AL_DFF_0 al_353f582f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[16]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[16]));
  AL_DFF_0 al_2dab617c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[17]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[17]));
  AL_DFF_0 al_cfbbadf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[44]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[44]));
  AL_DFF_0 al_2f21ee84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[45]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[45]));
  AL_DFF_0 al_7f9daeab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[46]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[46]));
  AL_DFF_0 al_ee2f6537 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b93da8d5[48]),
    .en(al_10206333[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dac85437[48]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    al_55ced1e7 (
    .a(al_28a9f919),
    .b(al_b93da8d5[0]),
    .c(al_53bb123b[0]),
    .d(al_3ee0d55a),
    .o(al_f11e0936));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    al_5a858798 (
    .a(al_28a9f919),
    .b(al_b93da8d5[1]),
    .c(al_53bb123b[1]),
    .d(al_3ee0d55a),
    .o(al_d017e8b1));
  AL_DFF_0 al_bbc15912 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f11e0936),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53bb123b[0]));
  AL_DFF_0 al_c47c188e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d017e8b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53bb123b[1]));
  AL_DFF_0 al_b27b1db8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_20b2d1cd[3]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_dd6ebfb0[3]));
  AL_DFF_0 al_25925e26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_20b2d1cd[4]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_dd6ebfb0[4]));
  AL_DFF_0 al_53a5afd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_20b2d1cd[0]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_dd6ebfb0[0]));
  AL_DFF_0 al_4a64930e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_20b2d1cd[1]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_dd6ebfb0[1]));
  AL_DFF_0 al_f8d36ede (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_20b2d1cd[2]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_dd6ebfb0[2]));
  AL_DFF_0 al_6653f298 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[11]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2602b5cf[3]));
  AL_DFF_0 al_91bf2c68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[12]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2602b5cf[4]));
  AL_DFF_0 al_e14e49d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[13]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2602b5cf[5]));
  AL_DFF_0 al_a133b58a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[14]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2602b5cf[6]));
  AL_DFF_0 al_bc489a30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[15]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2602b5cf[7]));
  AL_DFF_0 al_abf2ed95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[16]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2602b5cf[8]));
  AL_DFF_0 al_d12cee3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71f78ff1[17]),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_2602b5cf[9]));
  AL_DFF_0 al_a6df4eb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(rst),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c26eaf));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f3cffac0 (
    .i(al_a3c26eaf),
    .o(al_667181b3));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_37d2ed8b (
    .i(al_667181b3),
    .o(al_3ee0d55a));
  AL_DFF_0 al_22b2eab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4ecf439),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_456c110a));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*B*~(C)*D*E)"),
    .INIT(32'h0800fbcf))
    al_e0723559 (
    .a(al_cfaa4b74),
    .b(al_a67dc86a[0]),
    .c(al_a67dc86a[1]),
    .d(al_a67dc86a[2]),
    .e(al_81f91ff1[0]),
    .o(al_7711fc3[0]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haacaa0aa))
    al_9409fc0d (
    .a(al_4213cfc[4]),
    .b(al_2d60bf7c),
    .c(al_a67dc86a[0]),
    .d(al_a67dc86a[1]),
    .e(al_a67dc86a[2]),
    .o(al_7711fc3[4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_abf233bc (
    .a(al_7711fc3[4]),
    .b(al_7711fc3[3]),
    .c(al_7711fc3[2]),
    .d(al_7711fc3[1]),
    .e(al_7711fc3[0]),
    .o(al_96a13ff1));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~((F@E))+A*~(B)*~(C)*~(D)*~((F@E))+~(A)*B*~(C)*~(D)*~((F@E))+A*B*~(C)*~(D)*~((F@E))+~(A)*B*C*~(D)*~((F@E))+A*B*C*~(D)*~((F@E))+~(A)*~(B)*~(C)*D*~((F@E))+A*~(B)*~(C)*D*~((F@E))+A*B*~(C)*D*~((F@E))+~(A)*~(B)*C*D*~((F@E))+A*~(B)*C*D*~((F@E))+~(A)*B*C*D*~((F@E))+A*B*C*D*~((F@E))+A*B*~(C)*D*(F@E))"),
    .INIT(64'hfbcf08000800fbcf))
    al_e5341cf7 (
    .a(al_1c7e0f23),
    .b(al_a67dc86a[0]),
    .c(al_a67dc86a[1]),
    .d(al_a67dc86a[2]),
    .e(al_81f91ff1[0]),
    .f(al_81f91ff1[1]),
    .o(al_7711fc3[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C@(~B*~A))"),
    .INIT(8'h1e))
    al_5d98297f (
    .a(al_81f91ff1[0]),
    .b(al_81f91ff1[1]),
    .c(al_81f91ff1[2]),
    .o(al_edd1cf59));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55c55055))
    al_3cc15ad4 (
    .a(al_edd1cf59),
    .b(al_80cba1f),
    .c(al_a67dc86a[0]),
    .d(al_a67dc86a[1]),
    .e(al_a67dc86a[2]),
    .o(al_7711fc3[2]));
  AL_MAP_LUT4 #(
    .EQN("~(D@(~C*~B*~A))"),
    .INIT(16'h01fe))
    al_7f2fe4cb (
    .a(al_81f91ff1[0]),
    .b(al_81f91ff1[1]),
    .c(al_81f91ff1[2]),
    .d(al_81f91ff1[3]),
    .o(al_479ec121));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55c55055))
    al_215860f6 (
    .a(al_479ec121),
    .b(al_2f87218f),
    .c(al_a67dc86a[0]),
    .d(al_a67dc86a[1]),
    .e(al_a67dc86a[2]),
    .o(al_7711fc3[3]));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~C*~B*~A))"),
    .INIT(32'hfffe0001))
    al_9deeff24 (
    .a(al_81f91ff1[0]),
    .b(al_81f91ff1[1]),
    .c(al_81f91ff1[2]),
    .d(al_81f91ff1[3]),
    .e(al_81f91ff1[4]),
    .o(al_4213cfc[4]));
  AL_DFF_0 al_121cf1f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_96a13ff1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e620c305));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*A))"),
    .INIT(16'h007f))
    al_11f7b2e7 (
    .a(al_903070b1),
    .b(init_calib_complete),
    .c(al_90d84dc7[0]),
    .d(al_456c110a),
    .o(al_15b16fc6));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_9c887841 (
    .a(al_15b16fc6),
    .b(al_879aba03[0]),
    .o(al_e484293d[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*~A))"),
    .INIT(8'hb4))
    al_cf62691d (
    .a(al_15b16fc6),
    .b(al_879aba03[0]),
    .c(al_879aba03[1]),
    .o(al_e484293d[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_3546b89b (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_e484293d[0]),
    .d(al_e484293d[1]),
    .o(al_a4e4c65a));
  AL_DFF_0 al_4c42ca96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a4e4c65a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_df80405c));
  AL_DFF_0 al_9b3c8fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a9ec6721[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55b203da));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b4ed6e18 (
    .a(al_b4ecf439),
    .b(al_58fb4752[5]),
    .c(al_58851aab[0]),
    .o(al_3e489598[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_5dc494f5 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_146c01c2),
    .d(al_28de045),
    .e(al_7c3c9bb5),
    .f(al_24cee954),
    .o(al_6be20a95[0]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9e6375eb (
    .a(al_5453b759[1]),
    .b(al_3e489598[0]),
    .c(al_b9ba8b6c[0]),
    .o(al_28de045));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_87f45b01 (
    .a(al_5453b759[0]),
    .b(al_3e489598[0]),
    .c(al_77634075[0]),
    .o(al_146c01c2));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a0e9b70f (
    .a(al_5453b759[3]),
    .b(al_3e489598[0]),
    .c(al_d3350acc[0]),
    .o(al_7c3c9bb5));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_885d0222 (
    .a(al_3e489598[0]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[0]),
    .o(al_24cee954));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bba3aa71 (
    .a(al_b4ecf439),
    .b(al_58fb4752[6]),
    .c(al_58851aab[11]),
    .o(al_3e489598[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_a9c8aabd (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_bbfc232e),
    .d(al_3bb37542),
    .e(al_478a8b50),
    .f(al_de3eea8a),
    .o(al_6be20a95[11]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ddf5e034 (
    .a(al_5453b759[1]),
    .b(al_3e489598[11]),
    .c(al_b9ba8b6c[11]),
    .o(al_3bb37542));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_666c3255 (
    .a(al_5453b759[0]),
    .b(al_3e489598[11]),
    .c(al_77634075[11]),
    .o(al_bbfc232e));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b179b18d (
    .a(al_5453b759[3]),
    .b(al_3e489598[11]),
    .c(al_d3350acc[11]),
    .o(al_478a8b50));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_cbf1974c (
    .a(al_3e489598[11]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[11]),
    .o(al_de3eea8a));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9234b583 (
    .a(al_b4ecf439),
    .b(al_58fb4752[7]),
    .c(al_58851aab[12]),
    .o(al_3e489598[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_d2d3ff0c (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_1affa237),
    .d(al_77673c37),
    .e(al_30c9784a),
    .f(al_d253498d),
    .o(al_6be20a95[12]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_94593190 (
    .a(al_5453b759[1]),
    .b(al_3e489598[12]),
    .c(al_b9ba8b6c[12]),
    .o(al_77673c37));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_66448fb8 (
    .a(al_5453b759[0]),
    .b(al_3e489598[12]),
    .c(al_77634075[12]),
    .o(al_1affa237));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_56fcb2f8 (
    .a(al_5453b759[3]),
    .b(al_3e489598[12]),
    .c(al_d3350acc[12]),
    .o(al_30c9784a));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_1d97a3bf (
    .a(al_3e489598[12]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[12]),
    .o(al_d253498d));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c794d4d7 (
    .a(al_b4ecf439),
    .b(al_58fb4752[8]),
    .c(al_58851aab[13]),
    .o(al_3e489598[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_41a4ae8 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_63e01e1c),
    .d(al_15ef40b3),
    .e(al_e7da5efa),
    .f(al_4cd1569e),
    .o(al_6be20a95[13]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_8e072559 (
    .a(al_5453b759[1]),
    .b(al_3e489598[13]),
    .c(al_b9ba8b6c[13]),
    .o(al_15ef40b3));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_4f330ea2 (
    .a(al_5453b759[0]),
    .b(al_3e489598[13]),
    .c(al_77634075[13]),
    .o(al_63e01e1c));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_8cc946a5 (
    .a(al_5453b759[3]),
    .b(al_3e489598[13]),
    .c(al_d3350acc[13]),
    .o(al_e7da5efa));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_b4e90b8 (
    .a(al_3e489598[13]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[13]),
    .o(al_4cd1569e));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d902f2ca (
    .a(al_b4ecf439),
    .b(al_58fb4752[9]),
    .c(al_58851aab[14]),
    .o(al_3e489598[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_a3bb9216 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_8fe2ae6b),
    .d(al_8afb85c9),
    .e(al_1efa2be8),
    .f(al_5773cb6a),
    .o(al_6be20a95[14]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c7c83c97 (
    .a(al_5453b759[1]),
    .b(al_3e489598[14]),
    .c(al_b9ba8b6c[14]),
    .o(al_8afb85c9));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f1ff7489 (
    .a(al_5453b759[0]),
    .b(al_3e489598[14]),
    .c(al_77634075[14]),
    .o(al_8fe2ae6b));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_3e787214 (
    .a(al_5453b759[3]),
    .b(al_3e489598[14]),
    .c(al_d3350acc[14]),
    .o(al_1efa2be8));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_c25977e5 (
    .a(al_3e489598[14]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[14]),
    .o(al_5773cb6a));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_85fda17a (
    .a(al_b4ecf439),
    .b(al_58fb4752[10]),
    .c(al_58851aab[15]),
    .o(al_3e489598[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_2f2f94fd (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_1b24326b),
    .d(al_f589c903),
    .e(al_8fb41a59),
    .f(al_6ce9ade),
    .o(al_6be20a95[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_86fa233d (
    .a(al_5453b759[1]),
    .b(al_3e489598[15]),
    .c(al_b9ba8b6c[15]),
    .o(al_f589c903));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_553885ab (
    .a(al_5453b759[0]),
    .b(al_3e489598[15]),
    .c(al_77634075[15]),
    .o(al_1b24326b));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6469d939 (
    .a(al_5453b759[3]),
    .b(al_3e489598[15]),
    .c(al_d3350acc[15]),
    .o(al_8fb41a59));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_2da0d23a (
    .a(al_3e489598[15]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[15]),
    .o(al_6ce9ade));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_20ac0357 (
    .a(al_b4ecf439),
    .b(al_58fb4752[11]),
    .c(al_58851aab[16]),
    .o(al_3e489598[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_f2a546a6 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_4ba9f27d),
    .d(al_652e3f22),
    .e(al_693fd6e1),
    .f(al_8d59887e),
    .o(al_6be20a95[16]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_4f7bf1b1 (
    .a(al_5453b759[1]),
    .b(al_3e489598[16]),
    .c(al_b9ba8b6c[16]),
    .o(al_652e3f22));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_cd4167f6 (
    .a(al_5453b759[0]),
    .b(al_3e489598[16]),
    .c(al_77634075[16]),
    .o(al_4ba9f27d));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_71b12484 (
    .a(al_5453b759[3]),
    .b(al_3e489598[16]),
    .c(al_d3350acc[16]),
    .o(al_693fd6e1));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_83c0cb14 (
    .a(al_3e489598[16]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[16]),
    .o(al_8d59887e));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9020efee (
    .a(al_b4ecf439),
    .b(al_58fb4752[12]),
    .c(al_58851aab[17]),
    .o(al_3e489598[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_1b453b08 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_538ebf91),
    .d(al_cd9ec0c3),
    .e(al_2e98876c),
    .f(al_4417e3c3),
    .o(al_6be20a95[17]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d8bb362 (
    .a(al_5453b759[1]),
    .b(al_3e489598[17]),
    .c(al_b9ba8b6c[17]),
    .o(al_cd9ec0c3));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_51200744 (
    .a(al_5453b759[0]),
    .b(al_3e489598[17]),
    .c(al_77634075[17]),
    .o(al_538ebf91));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_34f258b1 (
    .a(al_5453b759[3]),
    .b(al_3e489598[17]),
    .c(al_d3350acc[17]),
    .o(al_2e98876c));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_3b54fb4c (
    .a(al_3e489598[17]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[17]),
    .o(al_4417e3c3));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_73d2468a (
    .a(al_b4ecf439),
    .b(al_58fb4752[3]),
    .c(al_58851aab[1]),
    .o(al_3e489598[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_3f4eaf1d (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_9fce8b6a),
    .d(al_6a20fb79),
    .e(al_7d8a45fd),
    .f(al_40c85aec),
    .o(al_6be20a95[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_44135179 (
    .a(al_5453b759[1]),
    .b(al_3e489598[1]),
    .c(al_b9ba8b6c[1]),
    .o(al_6a20fb79));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d3d1e2ba (
    .a(al_5453b759[0]),
    .b(al_3e489598[1]),
    .c(al_77634075[1]),
    .o(al_9fce8b6a));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c1d18b19 (
    .a(al_5453b759[3]),
    .b(al_3e489598[1]),
    .c(al_d3350acc[1]),
    .o(al_7d8a45fd));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_8f127b84 (
    .a(al_3e489598[1]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[1]),
    .o(al_40c85aec));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a3706b45 (
    .a(al_b4ecf439),
    .b(al_58fb4752[13]),
    .c(al_58851aab[24]),
    .o(al_3e489598[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_1cf4a545 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_3d802cc7),
    .d(al_751ac083),
    .e(al_fd225290),
    .f(al_f56597af),
    .o(al_6be20a95[24]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_65592e6c (
    .a(al_5453b759[1]),
    .b(al_3e489598[24]),
    .c(al_b9ba8b6c[24]),
    .o(al_751ac083));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e50e5830 (
    .a(al_5453b759[0]),
    .b(al_3e489598[24]),
    .c(al_77634075[24]),
    .o(al_3d802cc7));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6751705c (
    .a(al_5453b759[3]),
    .b(al_3e489598[24]),
    .c(al_d3350acc[24]),
    .o(al_fd225290));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_6edd9175 (
    .a(al_3e489598[24]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[24]),
    .o(al_f56597af));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_59b66b47 (
    .a(al_b4ecf439),
    .b(al_58fb4752[14]),
    .c(al_58851aab[25]),
    .o(al_3e489598[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_4e9de76d (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_10795ff8),
    .d(al_ac6abfed),
    .e(al_c45c98a0),
    .f(al_3fe6e16),
    .o(al_6be20a95[25]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e0e6807c (
    .a(al_5453b759[1]),
    .b(al_3e489598[25]),
    .c(al_b9ba8b6c[25]),
    .o(al_ac6abfed));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1b4ce45b (
    .a(al_5453b759[0]),
    .b(al_3e489598[25]),
    .c(al_77634075[25]),
    .o(al_10795ff8));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_63b813e3 (
    .a(al_5453b759[3]),
    .b(al_3e489598[25]),
    .c(al_d3350acc[25]),
    .o(al_c45c98a0));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_129a9c97 (
    .a(al_3e489598[25]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[25]),
    .o(al_3fe6e16));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_aba8d99b (
    .a(al_b4ecf439),
    .b(al_58fb4752[15]),
    .c(al_58851aab[26]),
    .o(al_3e489598[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_1a1245f6 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_fcdc6bd3),
    .d(al_c7d73a75),
    .e(al_92899c69),
    .f(al_3a54c9a1),
    .o(al_6be20a95[26]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d1884733 (
    .a(al_5453b759[1]),
    .b(al_3e489598[26]),
    .c(al_b9ba8b6c[26]),
    .o(al_c7d73a75));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f57959f (
    .a(al_5453b759[0]),
    .b(al_3e489598[26]),
    .c(al_77634075[26]),
    .o(al_fcdc6bd3));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6f65390b (
    .a(al_5453b759[3]),
    .b(al_3e489598[26]),
    .c(al_d3350acc[26]),
    .o(al_92899c69));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_1731c533 (
    .a(al_3e489598[26]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[26]),
    .o(al_3a54c9a1));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1c52483 (
    .a(al_b4ecf439),
    .b(al_58fb4752[16]),
    .c(al_58851aab[27]),
    .o(al_3e489598[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_f82b7874 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_3a2326ef),
    .d(al_3e34cef0),
    .e(al_f27a52ce),
    .f(al_b3f14729),
    .o(al_6be20a95[27]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_8d6f4b6d (
    .a(al_5453b759[1]),
    .b(al_3e489598[27]),
    .c(al_b9ba8b6c[27]),
    .o(al_3e34cef0));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_676c99d9 (
    .a(al_5453b759[0]),
    .b(al_3e489598[27]),
    .c(al_77634075[27]),
    .o(al_3a2326ef));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e76d3388 (
    .a(al_5453b759[3]),
    .b(al_3e489598[27]),
    .c(al_d3350acc[27]),
    .o(al_f27a52ce));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_12e89770 (
    .a(al_3e489598[27]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[27]),
    .o(al_b3f14729));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_106d104 (
    .a(al_b4ecf439),
    .b(al_58fb4752[17]),
    .c(al_58851aab[28]),
    .o(al_3e489598[28]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_ce89030 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_33769604),
    .d(al_44b901ea),
    .e(al_3ab8a708),
    .f(al_c83b5b3c),
    .o(al_6be20a95[28]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9263b974 (
    .a(al_5453b759[1]),
    .b(al_3e489598[28]),
    .c(al_b9ba8b6c[28]),
    .o(al_44b901ea));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ee146c3 (
    .a(al_5453b759[0]),
    .b(al_3e489598[28]),
    .c(al_77634075[28]),
    .o(al_33769604));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6c0d238a (
    .a(al_5453b759[3]),
    .b(al_3e489598[28]),
    .c(al_d3350acc[28]),
    .o(al_3ab8a708));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_debe1d1e (
    .a(al_3e489598[28]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[28]),
    .o(al_c83b5b3c));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_59c093c7 (
    .a(al_b4ecf439),
    .b(al_58fb4752[18]),
    .c(al_58851aab[29]),
    .o(al_3e489598[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_ac2ec647 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_616d30a),
    .d(al_bb4f41cb),
    .e(al_e20bf223),
    .f(al_70cc7b9e),
    .o(al_6be20a95[29]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c0168461 (
    .a(al_5453b759[1]),
    .b(al_3e489598[29]),
    .c(al_b9ba8b6c[29]),
    .o(al_bb4f41cb));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a98b4ae (
    .a(al_5453b759[0]),
    .b(al_3e489598[29]),
    .c(al_77634075[29]),
    .o(al_616d30a));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a34bbe3a (
    .a(al_5453b759[3]),
    .b(al_3e489598[29]),
    .c(al_d3350acc[29]),
    .o(al_e20bf223));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_ae897bef (
    .a(al_3e489598[29]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[29]),
    .o(al_70cc7b9e));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_23ae5a4b (
    .a(al_b4ecf439),
    .b(al_58fb4752[4]),
    .c(al_58851aab[2]),
    .o(al_3e489598[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_3c168680 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_6b420938),
    .d(al_fbff2df7),
    .e(al_f2acf56),
    .f(al_845e7508),
    .o(al_6be20a95[2]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b71fee9c (
    .a(al_5453b759[1]),
    .b(al_3e489598[2]),
    .c(al_b9ba8b6c[2]),
    .o(al_fbff2df7));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_af2a61c2 (
    .a(al_5453b759[0]),
    .b(al_3e489598[2]),
    .c(al_77634075[2]),
    .o(al_6b420938));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_763e6362 (
    .a(al_5453b759[3]),
    .b(al_3e489598[2]),
    .c(al_d3350acc[2]),
    .o(al_f2acf56));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_3b5fe982 (
    .a(al_3e489598[2]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[2]),
    .o(al_845e7508));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_546d6f59 (
    .a(al_b4ecf439),
    .b(al_58fb4752[19]),
    .c(al_58851aab[30]),
    .o(al_3e489598[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_7a377440 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_a9c6b32d),
    .d(al_799f406d),
    .e(al_445de8c8),
    .f(al_748564c9),
    .o(al_6be20a95[30]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9b066ad4 (
    .a(al_5453b759[1]),
    .b(al_3e489598[30]),
    .c(al_b9ba8b6c[30]),
    .o(al_799f406d));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_8a0c30f0 (
    .a(al_5453b759[0]),
    .b(al_3e489598[30]),
    .c(al_77634075[30]),
    .o(al_a9c6b32d));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_76e3983c (
    .a(al_5453b759[3]),
    .b(al_3e489598[30]),
    .c(al_d3350acc[30]),
    .o(al_445de8c8));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_de2f3257 (
    .a(al_3e489598[30]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[30]),
    .o(al_748564c9));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8536b34f (
    .a(al_b4ecf439),
    .b(al_58fb4752[20]),
    .c(al_58851aab[31]),
    .o(al_3e489598[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_d8af13a7 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_d66a1017),
    .d(al_95e1b9d1),
    .e(al_c304e63a),
    .f(al_8ad763a),
    .o(al_6be20a95[31]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_12af4696 (
    .a(al_5453b759[1]),
    .b(al_3e489598[31]),
    .c(al_b9ba8b6c[31]),
    .o(al_95e1b9d1));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ccb91709 (
    .a(al_5453b759[0]),
    .b(al_3e489598[31]),
    .c(al_77634075[31]),
    .o(al_d66a1017));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_dd60ddaa (
    .a(al_5453b759[3]),
    .b(al_3e489598[31]),
    .c(al_d3350acc[31]),
    .o(al_c304e63a));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_2bd06eb8 (
    .a(al_3e489598[31]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[31]),
    .o(al_8ad763a));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c4162bee (
    .a(al_b4ecf439),
    .b(al_58fb4752[21]),
    .c(al_58851aab[32]),
    .o(al_3e489598[32]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_529b7a4e (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_77bdc2db),
    .d(al_928fef0c),
    .e(al_38906f51),
    .f(al_ad0a7017),
    .o(al_6be20a95[32]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_70c76376 (
    .a(al_5453b759[1]),
    .b(al_3e489598[32]),
    .c(al_b9ba8b6c[32]),
    .o(al_928fef0c));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_5c0523c2 (
    .a(al_5453b759[0]),
    .b(al_3e489598[32]),
    .c(al_77634075[32]),
    .o(al_77bdc2db));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_5702095c (
    .a(al_5453b759[3]),
    .b(al_3e489598[32]),
    .c(al_d3350acc[32]),
    .o(al_38906f51));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_454b473e (
    .a(al_3e489598[32]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[32]),
    .o(al_ad0a7017));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ee332ed4 (
    .a(al_b4ecf439),
    .b(al_58fb4752[22]),
    .c(al_58851aab[33]),
    .o(al_3e489598[33]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_eff0fcfb (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_96a3d1d4),
    .d(al_445eda9d),
    .e(al_2770fee0),
    .f(al_5d634c36),
    .o(al_6be20a95[33]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a97e7af7 (
    .a(al_5453b759[1]),
    .b(al_3e489598[33]),
    .c(al_b9ba8b6c[33]),
    .o(al_445eda9d));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_69b3f41f (
    .a(al_5453b759[0]),
    .b(al_3e489598[33]),
    .c(al_77634075[33]),
    .o(al_96a3d1d4));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9449d978 (
    .a(al_5453b759[3]),
    .b(al_3e489598[33]),
    .c(al_d3350acc[33]),
    .o(al_2770fee0));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_ef5b126c (
    .a(al_3e489598[33]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[33]),
    .o(al_5d634c36));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e9ea7018 (
    .a(al_b4ecf439),
    .b(al_58fb4752[23]),
    .c(al_58851aab[34]),
    .o(al_3e489598[34]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_3e05c60 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_b6b5f546),
    .d(al_7f4f4920),
    .e(al_dac0f49d),
    .f(al_4f6e0352),
    .o(al_6be20a95[34]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_15017dc5 (
    .a(al_5453b759[1]),
    .b(al_3e489598[34]),
    .c(al_b9ba8b6c[34]),
    .o(al_7f4f4920));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_3b35dddc (
    .a(al_5453b759[0]),
    .b(al_3e489598[34]),
    .c(al_77634075[34]),
    .o(al_b6b5f546));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1c016ca5 (
    .a(al_5453b759[3]),
    .b(al_3e489598[34]),
    .c(al_d3350acc[34]),
    .o(al_dac0f49d));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_fd6e4148 (
    .a(al_3e489598[34]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[34]),
    .o(al_4f6e0352));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_615dc939 (
    .a(al_b4ecf439),
    .b(al_58fb4752[24]),
    .c(al_58851aab[35]),
    .o(al_3e489598[35]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_38ad0273 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_f15ca799),
    .d(al_374c386b),
    .e(al_e990f0b1),
    .f(al_49f2a7a7),
    .o(al_6be20a95[35]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_557accdf (
    .a(al_5453b759[1]),
    .b(al_3e489598[35]),
    .c(al_b9ba8b6c[35]),
    .o(al_374c386b));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_55d47232 (
    .a(al_5453b759[0]),
    .b(al_3e489598[35]),
    .c(al_77634075[35]),
    .o(al_f15ca799));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9666eb04 (
    .a(al_5453b759[3]),
    .b(al_3e489598[35]),
    .c(al_d3350acc[35]),
    .o(al_e990f0b1));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_9a6c4ae1 (
    .a(al_3e489598[35]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[35]),
    .o(al_49f2a7a7));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3ee6a4e (
    .a(al_b4ecf439),
    .b(al_58fb4752[25]),
    .c(al_58851aab[36]),
    .o(al_3e489598[36]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_842ff00 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_2c190380),
    .d(al_9906a30d),
    .e(al_3629f8f1),
    .f(al_a6dad665),
    .o(al_6be20a95[36]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_de982509 (
    .a(al_5453b759[1]),
    .b(al_3e489598[36]),
    .c(al_b9ba8b6c[36]),
    .o(al_9906a30d));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_8121c0ab (
    .a(al_5453b759[0]),
    .b(al_3e489598[36]),
    .c(al_77634075[36]),
    .o(al_2c190380));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ceb89b28 (
    .a(al_5453b759[3]),
    .b(al_3e489598[36]),
    .c(al_d3350acc[36]),
    .o(al_3629f8f1));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_c5ec8650 (
    .a(al_3e489598[36]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[36]),
    .o(al_a6dad665));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_49555af8 (
    .a(al_b4ecf439),
    .b(al_58fb4752[26]),
    .c(al_58851aab[37]),
    .o(al_3e489598[37]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_eee976f2 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_bc77e2de),
    .d(al_e089a5f3),
    .e(al_c9646708),
    .f(al_f6d87ba0),
    .o(al_6be20a95[37]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_80772487 (
    .a(al_5453b759[1]),
    .b(al_3e489598[37]),
    .c(al_b9ba8b6c[37]),
    .o(al_e089a5f3));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_27678a74 (
    .a(al_5453b759[0]),
    .b(al_3e489598[37]),
    .c(al_77634075[37]),
    .o(al_bc77e2de));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ecb1152a (
    .a(al_5453b759[3]),
    .b(al_3e489598[37]),
    .c(al_d3350acc[37]),
    .o(al_c9646708));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_224b450d (
    .a(al_3e489598[37]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[37]),
    .o(al_f6d87ba0));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_f19077a8 (
    .a(al_b4ecf439),
    .b(al_88a8db2c[0]),
    .o(al_3e489598[44]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_1efe8065 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_35747c43),
    .d(al_5f21f5b9),
    .e(al_d6220c5c),
    .f(al_90fdf0b2),
    .o(al_6be20a95[44]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c4f5ef2b (
    .a(al_5453b759[1]),
    .b(al_3e489598[44]),
    .c(al_b9ba8b6c[44]),
    .o(al_5f21f5b9));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a4af782f (
    .a(al_5453b759[0]),
    .b(al_3e489598[44]),
    .c(al_77634075[44]),
    .o(al_35747c43));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b7501341 (
    .a(al_5453b759[3]),
    .b(al_3e489598[44]),
    .c(al_d3350acc[44]),
    .o(al_d6220c5c));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_e1a49459 (
    .a(al_3e489598[44]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[44]),
    .o(al_90fdf0b2));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_556a4969 (
    .a(al_b4ecf439),
    .b(al_88a8db2c[1]),
    .o(al_3e489598[45]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_ae59c6b5 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_7bbf72a3),
    .d(al_f9c028af),
    .e(al_6969681f),
    .f(al_f6b9f88c),
    .o(al_6be20a95[45]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9e32cc43 (
    .a(al_5453b759[1]),
    .b(al_3e489598[45]),
    .c(al_b9ba8b6c[45]),
    .o(al_f9c028af));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b4f12334 (
    .a(al_5453b759[0]),
    .b(al_3e489598[45]),
    .c(al_77634075[45]),
    .o(al_7bbf72a3));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_62112e67 (
    .a(al_5453b759[3]),
    .b(al_3e489598[45]),
    .c(al_d3350acc[45]),
    .o(al_6969681f));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_1c367d18 (
    .a(al_3e489598[45]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[45]),
    .o(al_f6b9f88c));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_629adb2b (
    .a(al_b4ecf439),
    .b(al_88a8db2c[2]),
    .o(al_3e489598[46]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_1ad8c4e7 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_571561d4),
    .d(al_c0aba8fb),
    .e(al_1a076f81),
    .f(al_3fbbb328),
    .o(al_6be20a95[46]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c4fb43c2 (
    .a(al_5453b759[1]),
    .b(al_3e489598[46]),
    .c(al_b9ba8b6c[46]),
    .o(al_c0aba8fb));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9c398376 (
    .a(al_5453b759[0]),
    .b(al_3e489598[46]),
    .c(al_77634075[46]),
    .o(al_571561d4));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_271e88aa (
    .a(al_5453b759[3]),
    .b(al_3e489598[46]),
    .c(al_d3350acc[46]),
    .o(al_1a076f81));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_63deab5b (
    .a(al_3e489598[46]),
    .b(al_5453b759[2]),
    .c(al_9c434c4a[46]),
    .o(al_3fbbb328));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_beff6df7 (
    .a(al_49c007fc),
    .b(al_55b203da),
    .o(al_ff3a70dc));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b35d3f65 (
    .a(al_5453b759[3]),
    .b(al_b4ecf439),
    .c(al_d3350acc[48]),
    .o(al_10737a6f));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_65d2e4fd (
    .a(al_5453b759[2]),
    .b(al_b4ecf439),
    .c(al_9c434c4a[48]),
    .o(al_65b8bca5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h012389ab4567cdef))
    al_453fe987 (
    .a(al_765e8240[0]),
    .b(al_765e8240[1]),
    .c(al_84824ed8),
    .d(al_7546e20f),
    .e(al_10737a6f),
    .f(al_65b8bca5),
    .o(al_6be20a95[48]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_a528e160 (
    .a(al_ff3a70dc),
    .b(al_5c104e46),
    .o(al_b4ecf439));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_49cc4ae2 (
    .a(al_e484293d[0]),
    .b(al_879aba03[1]),
    .o(al_5453b759[3]));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*B*~(C)+A*~(B)*C)"),
    .INIT(8'h24))
    al_e0edd27b (
    .a(al_15b16fc6),
    .b(al_879aba03[0]),
    .c(al_879aba03[1]),
    .o(al_5453b759[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_c7d76ec6 (
    .a(al_e484293d[0]),
    .b(al_e484293d[1]),
    .o(al_5453b759[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_2554beba (
    .a(al_e484293d[0]),
    .b(al_879aba03[1]),
    .o(al_5453b759[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_65044bd2 (
    .a(al_5453b759[1]),
    .b(al_b4ecf439),
    .c(al_b9ba8b6c[48]),
    .o(al_7546e20f));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c03cb6b1 (
    .a(al_5453b759[0]),
    .b(al_b4ecf439),
    .c(al_77634075[48]),
    .o(al_84824ed8));
  AL_DFF_0 al_ec7333f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56e36fa5),
    .en(1'b1),
    .sr(al_3ee0d55a),
    .ss(1'b0),
    .q(al_bb796872));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_337be99a (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[0]),
    .d(al_4b620bb0[0]),
    .e(al_a5104c4f[0]),
    .f(al_dac85437[0]),
    .o(al_bbcf8fe1));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_5d4dff28 (
    .a(al_41ef913c),
    .b(al_457533f2),
    .c(al_e9f106ba),
    .d(al_bc420de3),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_3e1f1b94));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_d8c9ffd2 (
    .a(al_c952c11c),
    .b(al_e5cd290d),
    .c(al_1f4c68e6),
    .d(al_3c73e97d),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_a3d2c49d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_8a42f1a (
    .a(al_227f8a62),
    .b(al_c8afcceb),
    .c(al_e0aa83ea),
    .d(al_9f6af9ba),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_f7bf47b7));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_9b2f6fbe (
    .a(al_688aeb95),
    .b(al_bbfb7745),
    .c(al_b93da8d5[0]),
    .o(al_27d253fe));
  AL_MAP_LUT6 #(
    .EQN("(F@~(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'hf0cc55550f33aaaa))
    al_956c55a8 (
    .a(al_27d253fe),
    .b(al_1b8721f8),
    .c(al_b741880),
    .d(al_b93da8d5[0]),
    .e(al_b93da8d5[1]),
    .f(al_b93da8d5[24]),
    .o(al_57aea336));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_a0a4791a (
    .a(al_83d9c8d2),
    .b(al_232e33c9),
    .c(al_b93da8d5[0]),
    .o(al_e51d86f0));
  AL_MAP_LUT6 #(
    .EQN("(F@~(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'hf0cc55550f33aaaa))
    al_386e8afd (
    .a(al_e51d86f0),
    .b(al_95538c25),
    .c(al_b0e11bf3),
    .d(al_b93da8d5[0]),
    .e(al_b93da8d5[1]),
    .f(al_b93da8d5[35]),
    .o(al_7a27ca16));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_f74699fe (
    .a(al_a4dd8227),
    .b(al_97814ee2),
    .c(al_736e37f2),
    .d(al_f31ca00d),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_692dd432));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_1e5a3f74 (
    .a(al_ac3b1637),
    .b(al_f9500eb2),
    .c(al_9cb32c9b),
    .d(al_8ff2e306),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_dfa7ddb4));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_a82f614c (
    .a(al_4d37ff05),
    .b(al_50f5aee2),
    .c(al_c5c92715),
    .d(al_c7421999),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_4651c92a));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_df86d1ce (
    .a(al_bbcf8fe1),
    .b(al_8a415a42),
    .c(al_b93da8d5[0]),
    .o(al_71f78ff1[0]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_235cfb05 (
    .a(al_e769a1ac),
    .b(al_267ffb9b),
    .c(al_b93da8d5[0]),
    .o(al_504680b8));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_67526ee9 (
    .a(al_504680b8),
    .b(al_9e92954d),
    .c(al_bf6feeb3),
    .d(al_b93da8d5[0]),
    .e(al_b93da8d5[1]),
    .f(al_b93da8d5[26]),
    .o(al_7d5b642b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_2cd9f577 (
    .a(al_da2e6045),
    .b(al_2b60c4d7),
    .c(al_4f668848),
    .d(al_37cdc8a1),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_ebfbad28));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_8c93d5f1 (
    .a(al_533b1c82),
    .b(al_85770a25),
    .c(al_899fc7f2),
    .d(al_993b1b0f),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_98b1e60d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_ea194c55 (
    .a(al_ac45c87a),
    .b(al_2f21552f),
    .c(al_d17a0773),
    .d(al_3b11a186),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_8025a735));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_70003df5 (
    .a(al_8cae5877),
    .b(al_f71dba21),
    .c(al_b93da8d5[0]),
    .o(al_b681403c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_334a77cc (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[1]),
    .d(al_4b620bb0[1]),
    .e(al_a5104c4f[1]),
    .f(al_dac85437[1]),
    .o(al_2a1133de));
  AL_MAP_LUT6 #(
    .EQN("(F@~(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'hf0cc55550f33aaaa))
    al_11feba49 (
    .a(al_b681403c),
    .b(al_1f70c9fe),
    .c(al_d177c6b8),
    .d(al_b93da8d5[0]),
    .e(al_b93da8d5[1]),
    .f(al_b93da8d5[25]),
    .o(al_cc7cc536));
  AL_MAP_LUT6 #(
    .EQN("((F@C)*(E@B)*(D@A))"),
    .INIT(64'h0102040810204080))
    al_d2b6c12 (
    .a(al_3e1f1b94),
    .b(al_a3d2c49d),
    .c(al_4651c92a),
    .d(al_b93da8d5[31]),
    .e(al_b93da8d5[33]),
    .f(al_b93da8d5[37]),
    .o(al_e71d5665));
  AL_MAP_LUT6 #(
    .EQN("(B*A*(F@D)*(E@C))"),
    .INIT(64'h0008008008008000))
    al_96b24b32 (
    .a(al_7a27ca16),
    .b(al_cc7cc536),
    .c(al_ebfbad28),
    .d(al_98b1e60d),
    .e(al_b93da8d5[28]),
    .f(al_b93da8d5[30]),
    .o(al_93d3d349));
  AL_MAP_LUT6 #(
    .EQN("((E@C)*(F@B)*(D@A))"),
    .INIT(64'h0102102004084080))
    al_51c21dc (
    .a(al_3cb4c24d),
    .b(al_f7bf47b7),
    .c(al_8025a735),
    .d(al_b93da8d5[32]),
    .e(al_b93da8d5[34]),
    .f(al_b93da8d5[36]),
    .o(al_e54eae62));
  AL_MAP_LUT6 #(
    .EQN("(~B*A*(F@D)*(E@C))"),
    .INIT(64'h0002002002002000))
    al_f424393f (
    .a(al_57aea336),
    .b(al_7d5b642b),
    .c(al_692dd432),
    .d(al_dfa7ddb4),
    .e(al_b93da8d5[27]),
    .f(al_b93da8d5[29]),
    .o(al_b5b02afa));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_f3db4125 (
    .a(al_18326672),
    .b(al_5ec2c98e),
    .c(al_370aa1bb),
    .d(al_72b4a28e),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_ac74f6f1));
  AL_MAP_LUT6 #(
    .EQN("(~E*~A*~(F*~(D*C*B)))"),
    .INIT(64'h0000400000005555))
    al_b8a306ac (
    .a(al_ac74f6f1),
    .b(al_903070b1),
    .c(init_calib_complete),
    .d(al_90d84dc7[0]),
    .e(al_891340a1),
    .f(al_df80405c),
    .o(al_b6d031c2));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_3132a75d (
    .a(al_a67dc86a[0]),
    .b(al_a67dc86a[1]),
    .c(al_a67dc86a[2]),
    .o(al_718bc19f));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_d5659378 (
    .a(al_93d3d349),
    .b(al_b5b02afa),
    .c(al_e71d5665),
    .d(al_e54eae62),
    .e(al_b6d031c2),
    .f(al_718bc19f),
    .o(al_8bee4cd6));
  AL_MAP_LUT5 #(
    .EQN("~(C*~A*(~(B)*D*~(E)+B*~(D)*E+~(B)*D*E))"),
    .INIT(32'hefbfefff))
    al_263d977b (
    .a(al_891340a1),
    .b(al_a67dc86a[0]),
    .c(al_a67dc86a[1]),
    .d(al_a67dc86a[2]),
    .e(al_c360bf4c[0]),
    .o(al_954ec2c7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_52268c1c (
    .a(al_71f78ff1[0]),
    .b(al_71f78ff1[1]),
    .c(al_280c0ef0),
    .d(al_d2824414),
    .e(al_7cad9721),
    .f(al_681e3ff2),
    .o(al_4969cacc));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_c51ed175 (
    .a(al_2a1133de),
    .b(al_8a415a42),
    .c(al_b93da8d5[1]),
    .o(al_71f78ff1[1]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*~A))"),
    .INIT(16'h2333))
    al_505974e5 (
    .a(al_8bee4cd6),
    .b(al_4969cacc),
    .c(al_954ec2c7),
    .d(al_8a415a42),
    .o(al_74e913f6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_31bff99 (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[44]),
    .d(al_4b620bb0[44]),
    .e(al_a5104c4f[44]),
    .f(al_dac85437[44]),
    .o(al_895da8d));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_6e0a45ab (
    .a(al_895da8d),
    .b(al_8a415a42),
    .c(al_b93da8d5[44]),
    .o(al_da34749d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_3f68d89f (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[46]),
    .d(al_4b620bb0[46]),
    .e(al_a5104c4f[46]),
    .f(al_dac85437[46]),
    .o(al_1025128c));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_a271443e (
    .a(al_1025128c),
    .b(al_8a415a42),
    .c(al_b93da8d5[46]),
    .o(al_71f78ff1[46]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_6f8ee70a (
    .a(al_ffbe21a4[0]),
    .b(al_ffbe21a4[1]),
    .c(al_f0482f12[45]),
    .d(al_4b620bb0[45]),
    .e(al_a5104c4f[45]),
    .f(al_dac85437[45]),
    .o(al_691a84bb));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_9c823bfc (
    .a(al_61f44420),
    .b(ddr_app_rdy),
    .o(al_903070b1));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_3147cf88 (
    .a(al_691a84bb),
    .b(al_8a415a42),
    .c(al_b93da8d5[45]),
    .o(al_2d5968ed));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_cc2414dc (
    .a(al_da34749d),
    .b(al_71f78ff1[46]),
    .c(al_2d5968ed),
    .o(al_2bb5f88f));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_66962282 (
    .a(al_da34749d),
    .b(al_71f78ff1[46]),
    .c(al_2d5968ed),
    .d(al_c46598af[0]),
    .e(al_c46598af[1]),
    .o(al_8b4f323b));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~(C*~B*A)))"),
    .INIT(32'h00ff0020))
    al_45a2cabb (
    .a(al_74e913f6),
    .b(al_2bb5f88f),
    .c(al_8b4f323b),
    .d(al_1e3dbb5f),
    .e(al_bb796872),
    .o(al_56e36fa5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_c5420fc7 (
    .a(al_17bf017e),
    .b(al_5f86f74e),
    .c(al_fd00fe9e),
    .d(al_ece57492),
    .e(al_b93da8d5[0]),
    .f(al_b93da8d5[1]),
    .o(al_3cb4c24d));
  AL_DFF_0 al_b81c99ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b65fb56b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90d84dc7[1]));
  AL_DFF_0 al_4e2423bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aa1fb1d9),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_edb1c8b0));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_d8aa319d (
    .a(al_8ed48b41[0]),
    .b(al_8ed48b41[1]),
    .c(al_7a6f3e1[2]),
    .d(al_c6ae1e35[0]),
    .e(al_c6ae1e35[1]),
    .o(al_79fcd485[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_3001f645 (
    .a(al_48c3548d),
    .b(al_c360bf4c[1]),
    .o(al_aa1fb1d9));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(D*~(F@C)*~(E@B)))"),
    .INIT(64'h1555455551555455))
    al_af558c2b (
    .a(al_79fcd485[2]),
    .b(al_8ed48b41[0]),
    .c(al_8ed48b41[1]),
    .d(al_7a6f3e1[3]),
    .e(al_b56343fc[0]),
    .f(al_b56343fc[1]),
    .o(al_39c11c38));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_f9ff8ece (
    .a(al_8ed48b41[0]),
    .b(al_8ed48b41[1]),
    .c(al_7a6f3e1[1]),
    .d(al_393e4b3[0]),
    .e(al_393e4b3[1]),
    .o(al_79fcd485[1]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(D*~(F@C)*~(E@B)))"),
    .INIT(64'h1555455551555455))
    al_63b11d09 (
    .a(al_79fcd485[1]),
    .b(al_8ed48b41[0]),
    .c(al_8ed48b41[1]),
    .d(al_7a6f3e1[0]),
    .e(al_8664dd36[0]),
    .f(al_8664dd36[1]),
    .o(al_8a6a56f4));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E*~D))"),
    .INIT(32'h80008080))
    al_adbdc8a3 (
    .a(al_39c11c38),
    .b(al_8a6a56f4),
    .c(al_4db2fe90),
    .d(al_58d81d6c),
    .e(al_23659fe5),
    .o(al_856e8c85));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(~D*(A*C*~(E)*~(F)+A*C*~(E)*F+~(A)*~(C)*E*F+A*~(C)*E*F)))"),
    .INIT(64'h3330331333333313))
    al_42c318d5 (
    .a(al_856e8c85),
    .b(al_edb1c8b0),
    .c(al_c289c50a[0]),
    .d(al_c289c50a[1]),
    .e(al_c289c50a[2]),
    .f(al_ca5b8a7),
    .o(al_48c3548d));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*~A))"),
    .INIT(8'hc9))
    al_5fd3a27d (
    .a(al_6e677e24),
    .b(al_d712b15f),
    .c(al_1aabbc67),
    .o(al_cf086b44[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(~D*~B*~A))"),
    .INIT(16'hf0e1))
    al_29a69457 (
    .a(al_6e677e24),
    .b(al_d712b15f),
    .c(al_fd39d17d),
    .d(al_1aabbc67),
    .o(al_cf086b44[2]));
  AL_MAP_LUT6 #(
    .EQN("(E@(~F*~D*~C*~B*~A))"),
    .INIT(64'hffff0000fffe0001))
    al_77904c0b (
    .a(al_6e677e24),
    .b(al_d712b15f),
    .c(al_fd39d17d),
    .d(al_112c6aa0),
    .e(al_acf6f93e),
    .f(al_1aabbc67),
    .o(al_cf086b44[4]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_f3215200 (
    .a(al_6e677e24),
    .b(al_1aabbc67),
    .o(al_cf086b44[0]));
  AL_MAP_LUT5 #(
    .EQN("(D@(~E*~C*~B*~A))"),
    .INIT(32'hff00fe01))
    al_bc9ef1dc (
    .a(al_6e677e24),
    .b(al_d712b15f),
    .c(al_fd39d17d),
    .d(al_112c6aa0),
    .e(al_1aabbc67),
    .o(al_cf086b44[3]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_cda2e677 (
    .a(al_cf086b44[3]),
    .b(al_cf086b44[0]),
    .c(al_d712b15f),
    .d(al_fd39d17d),
    .e(al_acf6f93e),
    .o(al_dff56698[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_8dde4eb8 (
    .a(al_dff56698[0]),
    .b(al_1aabbc67),
    .o(al_886f442e[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_47847331 (
    .a(al_e42ac584[0]),
    .b(al_96dda245[0]),
    .c(al_535746d5[0]),
    .d(al_c8aa6814[0]),
    .e(al_40b9c486[0]),
    .f(al_40b9c486[1]),
    .o(al_b90e2b30[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_d9fc8b11 (
    .a(al_e42ac584[1]),
    .b(al_96dda245[1]),
    .c(al_535746d5[1]),
    .d(al_c8aa6814[1]),
    .e(al_40b9c486[0]),
    .f(al_40b9c486[1]),
    .o(al_b90e2b30[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_e11f4e2a (
    .a(al_e42ac584[2]),
    .b(al_96dda245[2]),
    .c(al_535746d5[2]),
    .d(al_c8aa6814[2]),
    .e(al_40b9c486[0]),
    .f(al_40b9c486[1]),
    .o(al_b90e2b30[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_2b9ee143 (
    .a(al_e42ac584[3]),
    .b(al_96dda245[3]),
    .c(al_535746d5[3]),
    .d(al_c8aa6814[3]),
    .e(al_40b9c486[0]),
    .f(al_40b9c486[1]),
    .o(al_b90e2b30[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_9a8c5acd (
    .a(al_e42ac584[4]),
    .b(al_96dda245[4]),
    .c(al_535746d5[4]),
    .d(al_c8aa6814[4]),
    .e(al_40b9c486[0]),
    .f(al_40b9c486[1]),
    .o(al_b90e2b30[4]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    al_84c36484 (
    .a(al_b4c6b3bd),
    .b(al_4a605a24[0]),
    .c(al_4a605a24[1]),
    .o(al_790e0f32));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_8186a789 (
    .a(al_790e0f32),
    .b(al_40b9c486[0]),
    .o(al_14c34e2f[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*~A))"),
    .INIT(8'hb4))
    al_7fd7f48c (
    .a(al_790e0f32),
    .b(al_40b9c486[0]),
    .c(al_40b9c486[1]),
    .o(al_14c34e2f[1]));
  AL_MAP_LUT4 #(
    .EQN("(D@(~C*~(B*~A)))"),
    .INIT(16'hf40b))
    al_40a9df2b (
    .a(al_75fd0159),
    .b(al_437081f2),
    .c(al_786dc891),
    .d(al_bd042336[0]),
    .o(al_bfcf9d28[0]));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~C*~(B*~A)))"),
    .INIT(32'hf4ff0b00))
    al_9b1e97bf (
    .a(al_75fd0159),
    .b(al_437081f2),
    .c(al_786dc891),
    .d(al_bd042336[0]),
    .e(al_bd042336[1]),
    .o(al_bfcf9d28[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_a1200bae (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_14c34e2f[0]),
    .d(al_14c34e2f[1]),
    .o(al_2057cd57));
  AL_DFF_0 al_fa79523 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2057cd57),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4c850aa));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(C*~A))"),
    .INIT(16'h639c))
    al_e7732776 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_14c34e2f[0]),
    .d(al_14c34e2f[1]),
    .o(al_89251c12[1]));
  AL_DFF_0 al_d559ff05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_89251c12[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25e1cc7));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_5fc0386e (
    .a(al_bd042336[0]),
    .b(al_bd042336[1]),
    .o(al_9119fd7[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(~E*~D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffffffcca0a0a080))
    al_c30fbf22 (
    .a(al_4396fcc1),
    .b(al_790e0f32),
    .c(al_9119fd7[0]),
    .d(al_40b9c486[0]),
    .e(al_40b9c486[1]),
    .f(al_7a6f3e1[0]),
    .o(al_c8d0e932[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_96acd1d0 (
    .a(al_bd042336[0]),
    .b(al_bd042336[1]),
    .o(al_9119fd7[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(~E*D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffffccffa0a080a0))
    al_415a8fec (
    .a(al_4396fcc1),
    .b(al_790e0f32),
    .c(al_9119fd7[1]),
    .d(al_40b9c486[0]),
    .e(al_40b9c486[1]),
    .f(al_7a6f3e1[1]),
    .o(al_c8d0e932[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6f14f189 (
    .a(al_bd042336[0]),
    .b(al_bd042336[1]),
    .o(al_9119fd7[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(E*~D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffccffffa080a0a0))
    al_814c85df (
    .a(al_4396fcc1),
    .b(al_790e0f32),
    .c(al_9119fd7[2]),
    .d(al_40b9c486[0]),
    .e(al_40b9c486[1]),
    .f(al_7a6f3e1[2]),
    .o(al_c8d0e932[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_a7b1a9cf (
    .a(al_bd042336[0]),
    .b(al_bd042336[1]),
    .o(al_9119fd7[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    al_e6f0111b (
    .a(al_75fd0159),
    .b(al_437081f2),
    .c(al_786dc891),
    .o(al_4396fcc1));
  AL_MAP_LUT6 #(
    .EQN("(~(E*D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hccffffff80a0a0a0))
    al_dbbf7b6b (
    .a(al_4396fcc1),
    .b(al_790e0f32),
    .c(al_9119fd7[3]),
    .d(al_40b9c486[0]),
    .e(al_40b9c486[1]),
    .f(al_7a6f3e1[3]),
    .o(al_c8d0e932[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_64dfc5ae (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[11]),
    .d(al_393e4b3[11]),
    .e(al_c6ae1e35[11]),
    .f(al_b56343fc[11]),
    .o(al_60f32aa5));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_c077b1ec (
    .a(al_60f32aa5),
    .b(al_e4c850aa),
    .c(al_8ed48b41[11]),
    .o(al_41f34c81[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_ab28d7c5 (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[12]),
    .d(al_393e4b3[12]),
    .e(al_c6ae1e35[12]),
    .f(al_b56343fc[12]),
    .o(al_d7c62deb));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_9c06fd09 (
    .a(al_d7c62deb),
    .b(al_e4c850aa),
    .c(al_8ed48b41[12]),
    .o(al_41f34c81[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_23f62d21 (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[13]),
    .d(al_393e4b3[13]),
    .e(al_c6ae1e35[13]),
    .f(al_b56343fc[13]),
    .o(al_53ec1776));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_bbdca306 (
    .a(al_53ec1776),
    .b(al_e4c850aa),
    .c(al_8ed48b41[13]),
    .o(al_41f34c81[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_dfd6554e (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[14]),
    .d(al_393e4b3[14]),
    .e(al_c6ae1e35[14]),
    .f(al_b56343fc[14]),
    .o(al_83399132));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_aad336f5 (
    .a(al_83399132),
    .b(al_e4c850aa),
    .c(al_8ed48b41[14]),
    .o(al_41f34c81[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_2aa0b7d3 (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[15]),
    .d(al_393e4b3[15]),
    .e(al_c6ae1e35[15]),
    .f(al_b56343fc[15]),
    .o(al_5aa41769));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_9d7360c6 (
    .a(al_5aa41769),
    .b(al_e4c850aa),
    .c(al_8ed48b41[15]),
    .o(al_41f34c81[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_51de68d9 (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[16]),
    .d(al_393e4b3[16]),
    .e(al_c6ae1e35[16]),
    .f(al_b56343fc[16]),
    .o(al_e69f53ab));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_7b59b3f (
    .a(al_e69f53ab),
    .b(al_e4c850aa),
    .c(al_8ed48b41[16]),
    .o(al_41f34c81[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_9bfa8c0b (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[17]),
    .d(al_393e4b3[17]),
    .e(al_c6ae1e35[17]),
    .f(al_b56343fc[17]),
    .o(al_86becd21));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_87866802 (
    .a(al_86becd21),
    .b(al_e4c850aa),
    .c(al_8ed48b41[17]),
    .o(al_41f34c81[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_11be002f (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[2]),
    .d(al_393e4b3[2]),
    .e(al_c6ae1e35[2]),
    .f(al_b56343fc[2]),
    .o(al_be3efaa4));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_1a52b366 (
    .a(al_be3efaa4),
    .b(al_e4c850aa),
    .c(al_8ed48b41[2]),
    .o(al_41f34c81[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_8afbf85e (
    .a(al_3b57d409[0]),
    .b(al_fc7c448b[0]),
    .c(al_d206e68[0]),
    .d(al_ce0a0d6b[0]),
    .e(al_66e5f5b5[0]),
    .f(al_66e5f5b5[1]),
    .o(al_100e6173));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_670c2587 (
    .a(al_100e6173),
    .b(al_58d81d6c),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[0]),
    .f(al_75c0d27f[0]),
    .o(al_c58f63f9[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_7a61c5e9 (
    .a(al_c58f63f9[0]),
    .b(al_fc7c448b[0]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_44b93047[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_98b9322a (
    .a(al_c58f63f9[0]),
    .b(al_ce0a0d6b[0]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_b6ac4cff[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_9fbdaaf0 (
    .a(al_c58f63f9[0]),
    .b(al_d206e68[0]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_4f585ca5[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_5109335e (
    .a(al_c58f63f9[0]),
    .b(al_3b57d409[0]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_526d80ee[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_4db1f027 (
    .a(al_44b93047[0]),
    .b(al_b6ac4cff[0]),
    .c(al_4f585ca5[0]),
    .d(al_526d80ee[0]),
    .e(al_bd042336[0]),
    .f(al_bd042336[1]),
    .o(al_8023991e[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_72edb4a1 (
    .a(al_3b57d409[1]),
    .b(al_fc7c448b[1]),
    .c(al_d206e68[1]),
    .d(al_ce0a0d6b[1]),
    .e(al_66e5f5b5[0]),
    .f(al_66e5f5b5[1]),
    .o(al_1a4dce1b));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_b4be9906 (
    .a(al_1a4dce1b),
    .b(al_58d81d6c),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[1]),
    .f(al_75c0d27f[1]),
    .o(al_c58f63f9[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_bdbe2fa3 (
    .a(al_c58f63f9[1]),
    .b(al_fc7c448b[1]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_44b93047[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_1670ae (
    .a(al_c58f63f9[1]),
    .b(al_ce0a0d6b[1]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_b6ac4cff[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_dadda443 (
    .a(al_c58f63f9[1]),
    .b(al_d206e68[1]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_4f585ca5[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_343965cd (
    .a(al_c58f63f9[1]),
    .b(al_3b57d409[1]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_526d80ee[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_5976d41a (
    .a(al_44b93047[1]),
    .b(al_b6ac4cff[1]),
    .c(al_4f585ca5[1]),
    .d(al_526d80ee[1]),
    .e(al_bd042336[0]),
    .f(al_bd042336[1]),
    .o(al_8023991e[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_c3b8de5b (
    .a(al_3b57d409[2]),
    .b(al_fc7c448b[2]),
    .c(al_d206e68[2]),
    .d(al_ce0a0d6b[2]),
    .e(al_66e5f5b5[0]),
    .f(al_66e5f5b5[1]),
    .o(al_b0d45bcf));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_86c71c80 (
    .a(al_b0d45bcf),
    .b(al_58d81d6c),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[2]),
    .f(al_75c0d27f[2]),
    .o(al_c58f63f9[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_8456011 (
    .a(al_c58f63f9[2]),
    .b(al_fc7c448b[2]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_44b93047[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_74ed580c (
    .a(al_c58f63f9[2]),
    .b(al_ce0a0d6b[2]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_b6ac4cff[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_fa102d1d (
    .a(al_c58f63f9[2]),
    .b(al_d206e68[2]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_4f585ca5[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_e664382e (
    .a(al_c58f63f9[2]),
    .b(al_3b57d409[2]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_526d80ee[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_2e329344 (
    .a(al_44b93047[2]),
    .b(al_b6ac4cff[2]),
    .c(al_4f585ca5[2]),
    .d(al_526d80ee[2]),
    .e(al_bd042336[0]),
    .f(al_bd042336[1]),
    .o(al_8023991e[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_3aa5d3a5 (
    .a(al_3b57d409[3]),
    .b(al_fc7c448b[3]),
    .c(al_d206e68[3]),
    .d(al_ce0a0d6b[3]),
    .e(al_66e5f5b5[0]),
    .f(al_66e5f5b5[1]),
    .o(al_b13009b2));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_f5202888 (
    .a(al_b13009b2),
    .b(al_58d81d6c),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[3]),
    .f(al_75c0d27f[3]),
    .o(al_c58f63f9[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_99b3a4e9 (
    .a(al_c58f63f9[3]),
    .b(al_fc7c448b[3]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_44b93047[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_4e7ecf1b (
    .a(al_c58f63f9[3]),
    .b(al_ce0a0d6b[3]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_b6ac4cff[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_a3059340 (
    .a(al_c58f63f9[3]),
    .b(al_d206e68[3]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_4f585ca5[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_32b07030 (
    .a(al_c58f63f9[3]),
    .b(al_3b57d409[3]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_526d80ee[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_f6e02777 (
    .a(al_44b93047[3]),
    .b(al_b6ac4cff[3]),
    .c(al_4f585ca5[3]),
    .d(al_526d80ee[3]),
    .e(al_bd042336[0]),
    .f(al_bd042336[1]),
    .o(al_8023991e[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_1a4c42e4 (
    .a(al_3b57d409[4]),
    .b(al_fc7c448b[4]),
    .c(al_d206e68[4]),
    .d(al_ce0a0d6b[4]),
    .e(al_66e5f5b5[0]),
    .f(al_66e5f5b5[1]),
    .o(al_aecd56b));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*(D@C)))*~(B)+~A*(E*(D@C))*~(B)+~(~A)*(E*(D@C))*B+~A*(E*(D@C))*B)"),
    .INIT(32'h1dd11111))
    al_e385fb0b (
    .a(al_aecd56b),
    .b(al_58d81d6c),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[4]),
    .o(al_c58f63f9[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_5808d1fe (
    .a(al_c58f63f9[4]),
    .b(al_fc7c448b[4]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_44b93047[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_52d30158 (
    .a(al_c58f63f9[4]),
    .b(al_ce0a0d6b[4]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_b6ac4cff[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_c4cc0f56 (
    .a(al_c58f63f9[4]),
    .b(al_d206e68[4]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_4f585ca5[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_c2d4f7e3 (
    .a(al_c58f63f9[4]),
    .b(al_3b57d409[4]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_526d80ee[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_391ee9f4 (
    .a(al_44b93047[4]),
    .b(al_b6ac4cff[4]),
    .c(al_4f585ca5[4]),
    .d(al_526d80ee[4]),
    .e(al_bd042336[0]),
    .f(al_bd042336[1]),
    .o(al_8023991e[4]));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*A*~(E*~D))"),
    .INIT(32'h08000808))
    al_518fb65f (
    .a(al_39c11c38),
    .b(al_8a6a56f4),
    .c(al_4db2fe90),
    .d(al_58d81d6c),
    .e(al_23659fe5),
    .o(al_128dcf82));
  AL_MAP_LUT6 #(
    .EQN("(F*~(E*D*C*B*A))"),
    .INIT(64'h7fffffff00000000))
    al_69b4c817 (
    .a(al_8d6dd847),
    .b(al_f22292ec),
    .c(al_6f281a7f),
    .d(al_d94dff22),
    .e(al_ef2f822e),
    .f(al_c289c50a[0]),
    .o(al_c7a5b233));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*B*~(E*A)))"),
    .INIT(32'h00bf003f))
    al_3f4abbde (
    .a(al_25e1cc7),
    .b(al_c289c50a[0]),
    .c(al_c289c50a[1]),
    .d(al_c289c50a[2]),
    .e(al_c360bf4c[1]),
    .o(al_79fd4e7c));
  AL_MAP_LUT6 #(
    .EQN("(~D*~(F*~(~E*~(C*~(~B*~A)))))"),
    .INIT(64'h0000001f00ff00ff))
    al_b242342d (
    .a(al_5b931dce),
    .b(al_8f446276),
    .c(al_c7a5b233),
    .d(al_7393f55f),
    .e(al_5ab672a4),
    .f(al_79fd4e7c),
    .o(al_57cd6e45[0]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*D*C*B))"),
    .INIT(32'h2aaaaaaa))
    al_24350fbb (
    .a(al_128dcf82),
    .b(al_8d6dd847),
    .c(al_f22292ec),
    .d(al_6f281a7f),
    .e(al_d94dff22),
    .o(al_5b931dce));
  AL_MAP_LUT4 #(
    .EQN("(A*(~(B)*~(C)*~(D)+B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D+~(B)*C*D))"),
    .INIT(16'h282a))
    al_df6b83f5 (
    .a(al_786dc891),
    .b(al_c289c50a[0]),
    .c(al_c289c50a[1]),
    .d(al_ca5b8a7),
    .o(al_7393f55f));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~(~D*~(C*~(F*~(~B*A)))))"),
    .INIT(64'hffff00dfffff000f))
    al_a898a882 (
    .a(al_58fb4752[3]),
    .b(al_58fb4752[4]),
    .c(al_f7a41bbb),
    .d(al_c289c50a[0]),
    .e(al_c289c50a[1]),
    .f(al_23659fe5),
    .o(al_5ab672a4));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_e35a89b7 (
    .a(al_856e8c85),
    .b(al_6896ad14),
    .c(al_23659fe5),
    .o(al_8f446276));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~A))*~(B)+D*(C*~A)*~(B)+~(D)*(C*~A)*B+D*(C*~A)*B)"),
    .INIT(16'h7340))
    al_b6f218d8 (
    .a(al_25e1cc7),
    .b(al_c289c50a[0]),
    .c(al_c360bf4c[1]),
    .d(al_8932a489),
    .o(al_cd0e3f19));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h03f0aaff03ffaaff))
    al_2340764e (
    .a(al_cd0e3f19),
    .b(al_25e1cc7),
    .c(al_c289c50a[0]),
    .d(al_c289c50a[1]),
    .e(al_c289c50a[2]),
    .f(al_ca5b8a7),
    .o(al_2e2c5e0e));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(~E*D*~(~B*~A)))"),
    .INIT(32'h0f0fef0f))
    al_761f3221 (
    .a(al_5b931dce),
    .b(al_856e8c85),
    .c(al_2e2c5e0e),
    .d(al_fbe54a4d),
    .e(al_c289c50a[2]),
    .o(al_57cd6e45[1]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    al_a1a1a8d5 (
    .a(al_25e1cc7),
    .b(al_c289c50a[0]),
    .c(al_c360bf4c[1]),
    .d(al_8932a489),
    .o(al_161ea611));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfcf05500fcff5500))
    al_2775824f (
    .a(al_161ea611),
    .b(al_25e1cc7),
    .c(al_c289c50a[0]),
    .d(al_c289c50a[1]),
    .e(al_c289c50a[2]),
    .f(al_ca5b8a7),
    .o(al_57cd6e45[2]));
  AL_MAP_LUT5 #(
    .EQN("((~B*A)*~(C)*~(D)*~(E)+(~B*A)*C*~(D)*~(E)+~((~B*A))*~(C)*D*~(E)+(~B*A)*~(C)*D*~(E)+~((~B*A))*C*~(D)*E+(~B*A)*C*~(D)*E+~((~B*A))*~(C)*D*E+(~B*A)*~(C)*D*E+~((~B*A))*C*D*E+(~B*A)*C*D*E)"),
    .INIT(32'hfff00f22))
    al_75ce1b3c (
    .a(al_c20a9a7e),
    .b(al_56be2a2c),
    .c(al_b4c6b3bd),
    .d(al_4a605a24[0]),
    .e(al_4a605a24[1]),
    .o(al_90c83bf9[0]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(~C*B*A))"),
    .INIT(16'hff08))
    al_fc49e80d (
    .a(al_c20a9a7e),
    .b(al_56be2a2c),
    .c(al_4a605a24[0]),
    .d(al_4a605a24[1]),
    .o(al_90c83bf9[1]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_bf07e9c1 (
    .a(al_ee675012),
    .b(al_d2b50474),
    .c(al_38fc89af),
    .o(al_9cbe46a));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_8d3c6d6a (
    .a(al_681de671),
    .b(al_d2b50474),
    .c(al_38fc89af),
    .o(al_9ccb16fd));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_bca7f114 (
    .a(al_6d851644),
    .b(al_d2b50474),
    .c(al_38fc89af),
    .o(al_da6c82d));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_4afb44bd (
    .a(al_cf11b78b[1]),
    .b(al_c289c50a[0]),
    .c(al_c289c50a[1]),
    .d(al_c289c50a[2]),
    .e(al_898823b1),
    .o(al_d2b50474));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_72145f5f (
    .a(al_5b2f4c49),
    .b(al_d2b50474),
    .c(al_38fc89af),
    .o(al_f68c5dd8));
  AL_DFF_0 al_8d8af24f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6237c511),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_ef9d2d1b));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    al_a6bf542a (
    .a(al_10f0cebf),
    .b(al_ef9d2d1b),
    .c(al_8932a489),
    .o(al_6237c511));
  AL_DFF_0 al_af42ced2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf086b44[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_6e677e24));
  AL_DFF_0 al_ad788bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf086b44[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_d712b15f));
  AL_DFF_0 al_3d413503 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf086b44[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_fd39d17d));
  AL_DFF_0 al_250fb452 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf086b44[3]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_112c6aa0));
  AL_DFF_0 al_75f524e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf086b44[4]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_acf6f93e));
  AL_DFF_0 al_999d855 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a119035a[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7f004572));
  AL_DFF_0 al_f231a37e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a119035a[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1827053f));
  AL_DFF_0 al_80aa6b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a119035a[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2934d890));
  AL_DFF_0 al_98998d06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a119035a[3]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_3d0b7065));
  AL_DFF_0 al_783011ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_640bf3cc[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_176b7b0e));
  AL_DFF_0 al_4cddaafd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_640bf3cc[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7c2107c8));
  AL_DFF_0 al_f632dab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_640bf3cc[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_5f82f20d));
  AL_DFF_0 al_ac47601b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_640bf3cc[3]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_dd0180f1));
  AL_DFF_0 al_6d45d765 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3cc6453[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_947ff24d));
  AL_DFF_0 al_9b05d32e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3cc6453[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_816f1763));
  AL_DFF_0 al_f201d83f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3cc6453[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_d840d9f3));
  AL_DFF_0 al_cedb4042 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3cc6453[3]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_38e5040b));
  AL_DFF_0 al_b6e13210 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_259bb519[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2b09146));
  AL_DFF_0 al_2e9e52b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_259bb519[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_eba4eddb));
  AL_DFF_0 al_873c5e9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_259bb519[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_55cda68f));
  AL_DFF_0 al_f631b4f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_259bb519[3]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_e7ff6740));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_48856bc7 (
    .a(al_c289c50a[0]),
    .b(al_c289c50a[1]),
    .c(al_c289c50a[2]),
    .o(al_4c28a161));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_c625eb82 (
    .a(al_4c28a161),
    .b(al_8ed48b41[0]),
    .c(al_8ed48b41[1]),
    .o(al_681de671));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5fd361a9 (
    .a(al_681de671),
    .b(al_c360bf4c[1]),
    .o(al_ff84082));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_7fb9ce87 (
    .a(al_ff84082),
    .b(al_176b7b0e),
    .c(al_7c2107c8),
    .d(al_5f82f20d),
    .e(al_dd0180f1),
    .f(al_3fdd9bd4),
    .o(al_640bf3cc[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_9c4da3bd (
    .a(al_ff84082),
    .b(al_176b7b0e),
    .c(al_3fdd9bd4),
    .o(al_640bf3cc[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_810dd008 (
    .a(al_ff84082),
    .b(al_176b7b0e),
    .c(al_7c2107c8),
    .d(al_3fdd9bd4),
    .o(al_640bf3cc[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_552fd80e (
    .a(al_ff84082),
    .b(al_176b7b0e),
    .c(al_7c2107c8),
    .d(al_5f82f20d),
    .e(al_3fdd9bd4),
    .o(al_640bf3cc[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_1e9f78f8 (
    .a(al_4c28a161),
    .b(al_8ed48b41[0]),
    .c(al_8ed48b41[1]),
    .o(al_6d851644));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_dcf1712 (
    .a(al_6d851644),
    .b(al_c360bf4c[1]),
    .o(al_49045baf));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_c03bd66d (
    .a(al_49045baf),
    .b(al_947ff24d),
    .c(al_816f1763),
    .d(al_d840d9f3),
    .e(al_38e5040b),
    .f(al_724e96cb),
    .o(al_c3cc6453[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_53d05f19 (
    .a(al_49045baf),
    .b(al_947ff24d),
    .c(al_724e96cb),
    .o(al_c3cc6453[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_8132ffc9 (
    .a(al_49045baf),
    .b(al_947ff24d),
    .c(al_816f1763),
    .d(al_724e96cb),
    .o(al_c3cc6453[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_6d8671ba (
    .a(al_49045baf),
    .b(al_947ff24d),
    .c(al_816f1763),
    .d(al_d840d9f3),
    .e(al_724e96cb),
    .o(al_c3cc6453[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_812ead21 (
    .a(al_4c28a161),
    .b(al_8ed48b41[0]),
    .c(al_8ed48b41[1]),
    .o(al_5b2f4c49));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_3a5b9020 (
    .a(al_5b2f4c49),
    .b(al_c360bf4c[1]),
    .o(al_43b9e423));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_96ce80ae (
    .a(al_43b9e423),
    .b(al_2b09146),
    .c(al_eba4eddb),
    .d(al_55cda68f),
    .e(al_e7ff6740),
    .f(al_f6cbc027),
    .o(al_259bb519[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_215f7c6a (
    .a(al_43b9e423),
    .b(al_2b09146),
    .c(al_f6cbc027),
    .o(al_259bb519[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_96dd8055 (
    .a(al_43b9e423),
    .b(al_2b09146),
    .c(al_eba4eddb),
    .d(al_f6cbc027),
    .o(al_259bb519[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_f9fa61af (
    .a(al_43b9e423),
    .b(al_2b09146),
    .c(al_eba4eddb),
    .d(al_55cda68f),
    .e(al_f6cbc027),
    .o(al_259bb519[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_84f4508 (
    .a(al_4c28a161),
    .b(al_8ed48b41[0]),
    .c(al_8ed48b41[1]),
    .o(al_ee675012));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_c40c8278 (
    .a(al_ee675012),
    .b(al_c360bf4c[1]),
    .o(al_7a822c74));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_b8bcf17b (
    .a(al_7a822c74),
    .b(al_7f004572),
    .c(al_1827053f),
    .d(al_2934d890),
    .e(al_3d0b7065),
    .f(al_51ceabf0),
    .o(al_a119035a[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_cc73bf4f (
    .a(al_7a822c74),
    .b(al_7f004572),
    .c(al_51ceabf0),
    .o(al_a119035a[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_9e5d6465 (
    .a(al_7a822c74),
    .b(al_7f004572),
    .c(al_1827053f),
    .d(al_51ceabf0),
    .o(al_a119035a[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_fc58937e (
    .a(al_7a822c74),
    .b(al_7f004572),
    .c(al_1827053f),
    .d(al_2934d890),
    .e(al_51ceabf0),
    .o(al_a119035a[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_4e5d8e89 (
    .a(al_640bf3cc[3]),
    .b(al_640bf3cc[0]),
    .c(al_640bf3cc[1]),
    .d(al_640bf3cc[2]),
    .o(al_8a6bb27f[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_a0ed9a61 (
    .a(al_c3cc6453[3]),
    .b(al_c3cc6453[0]),
    .c(al_c3cc6453[1]),
    .d(al_c3cc6453[2]),
    .o(al_8a6bb27f[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_b4d063e1 (
    .a(al_259bb519[3]),
    .b(al_259bb519[0]),
    .c(al_259bb519[1]),
    .d(al_259bb519[2]),
    .o(al_8a6bb27f[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_9775559d (
    .a(al_a119035a[3]),
    .b(al_a119035a[0]),
    .c(al_a119035a[1]),
    .d(al_a119035a[2]),
    .o(al_8a6bb27f[0]));
  AL_DFF_0 al_a590fc79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8a6bb27f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51ceabf0));
  AL_DFF_0 al_f8e0cb7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8a6bb27f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3fdd9bd4));
  AL_DFF_0 al_c93a0236 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8a6bb27f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_724e96cb));
  AL_DFF_0 al_b00cb392 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8a6bb27f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f6cbc027));
  AL_DFF_0 al_efac456d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a3d2fd0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56598d));
  AL_DFF_0 al_d784b727 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[24]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_868dabaf));
  AL_DFF_0 al_45d56675 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[25]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_46fc25e7));
  AL_DFF_0 al_26c22a5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[26]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_22d551b1));
  AL_DFF_0 al_1888b097 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[27]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_af3a3adf));
  AL_DFF_0 al_b2a940be (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[28]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_80336d41));
  AL_DFF_0 al_d0fe3695 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[29]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_fe185597));
  AL_DFF_0 al_c46172e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[30]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_cf63226f));
  AL_DFF_0 al_57aa6ee0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[31]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_88d2570b));
  AL_DFF_0 al_e1ebdf7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[32]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1ea50fd5));
  AL_DFF_0 al_a9600593 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[33]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_cf05798c));
  AL_DFF_0 al_af17d033 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[34]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_627e01b));
  AL_DFF_0 al_397f2a1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[35]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9a04ce8f));
  AL_DFF_0 al_849b88a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[36]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7aadf07));
  AL_DFF_0 al_43bdff77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[37]),
    .en(al_9cbe46a),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_ab1b96f9));
  AL_DFF_0 al_74d338c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f8a12fba),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_122466dd));
  AL_DFF_0 al_d5775257 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[24]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_25fc271e));
  AL_DFF_0 al_15d4f1c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[25]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_fb20038d));
  AL_DFF_0 al_8398e186 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[26]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_ffaa6ed4));
  AL_DFF_0 al_16ebef00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[27]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9384d2a6));
  AL_DFF_0 al_c0838b90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[28]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_5bb79c4f));
  AL_DFF_0 al_9722f865 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[29]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_f0cf2c1b));
  AL_DFF_0 al_c11735fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[30]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_a0f44394));
  AL_DFF_0 al_86d2bb62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[31]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_ae9de7f7));
  AL_DFF_0 al_65433635 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[32]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_48347124));
  AL_DFF_0 al_bf99563b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[33]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_ddc7a73f));
  AL_DFF_0 al_5019ec9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[34]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_58f4bcca));
  AL_DFF_0 al_2b3a1def (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[35]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_4c783ffb));
  AL_DFF_0 al_af5d612a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[36]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_b7e2e71f));
  AL_DFF_0 al_f0048341 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[37]),
    .en(al_9ccb16fd),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_c34f057a));
  AL_DFF_0 al_a17abc6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_45523d4b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_195fd12));
  AL_DFF_0 al_bd049cde (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[24]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_81d476eb));
  AL_DFF_0 al_6f6c8ae2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[25]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f586c30));
  AL_DFF_0 al_53b6a3ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[26]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_f53cd64f));
  AL_DFF_0 al_4fcc96ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[27]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_5c212f53));
  AL_DFF_0 al_56107ef1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[28]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_b6b9db4));
  AL_DFF_0 al_b6a0de0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[29]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_b797198c));
  AL_DFF_0 al_dbfb13d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[30]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_73f87281));
  AL_DFF_0 al_597f3a96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[31]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_cafe0ec3));
  AL_DFF_0 al_82150122 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[32]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_67f78c15));
  AL_DFF_0 al_d34f17a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[33]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_a620188b));
  AL_DFF_0 al_7284d00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[34]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_a5fb3197));
  AL_DFF_0 al_22e6485d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[35]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_38c33a99));
  AL_DFF_0 al_b4207094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[36]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_5cd3a57d));
  AL_DFF_0 al_9122dc97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[37]),
    .en(al_da6c82d),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_fccfd8ff));
  AL_DFF_0 al_7a717c63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_451ab1e2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_91e55879));
  AL_DFF_0 al_f430ebd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[24]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_699f3bb8));
  AL_DFF_0 al_88d76a80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[25]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_4ce39135));
  AL_DFF_0 al_c9884697 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[26]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_b93ffb04));
  AL_DFF_0 al_ec383053 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[27]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_d8c260df));
  AL_DFF_0 al_1ccbbd98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[28]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_42cfbe9b));
  AL_DFF_0 al_3705e8a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[29]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_8b71d8b7));
  AL_DFF_0 al_ed909e53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[30]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_79ca7989));
  AL_DFF_0 al_bc371409 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[31]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_3c683e0a));
  AL_DFF_0 al_38988e2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[32]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_3b14a515));
  AL_DFF_0 al_2cac7dbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[33]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_79ced939));
  AL_DFF_0 al_2e47fe51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[34]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_865e3224));
  AL_DFF_0 al_198a7163 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[35]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_310a635));
  AL_DFF_0 al_7e48b613 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[36]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_b2200d60));
  AL_DFF_0 al_ed91ffe6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[37]),
    .en(al_f68c5dd8),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_be66ece6));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_d435cb2f (
    .a(al_681de671),
    .b(al_d2b50474),
    .c(al_122466dd),
    .d(al_38fc89af),
    .e(al_18fc9355),
    .o(al_f8a12fba));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_cb10a3d4 (
    .a(al_ee675012),
    .b(al_d2b50474),
    .c(al_b56598d),
    .d(al_38fc89af),
    .e(al_18fc9355),
    .o(al_1a3d2fd0));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_f0e4c7ba (
    .a(al_5b2f4c49),
    .b(al_d2b50474),
    .c(al_91e55879),
    .d(al_38fc89af),
    .e(al_18fc9355),
    .o(al_451ab1e2));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_824da15a (
    .a(al_6d851644),
    .b(al_d2b50474),
    .c(al_195fd12),
    .d(al_38fc89af),
    .e(al_18fc9355),
    .o(al_45523d4b));
  AL_DFF_0 al_c8516d46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_886f442e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_38fc89af));
  AL_DFF_0 al_25bcec9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dff56698[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1aabbc67));
  AL_DFF_0 al_6fb60a90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dfc7aeab),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_d50c8b50));
  AL_MAP_LUT6 #(
    .EQN("(~C*~(~D*~(~F*~E*B*A)))"),
    .INIT(64'h0f000f000f000f08))
    al_3bf960d1 (
    .a(al_c20a9a7e),
    .b(al_cd0bc85d),
    .c(al_b4c6b3bd),
    .d(al_d50c8b50),
    .e(al_4a605a24[0]),
    .f(al_4a605a24[1]),
    .o(al_dfc7aeab));
  AL_DFF_0 al_4271b987 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ce5f7b78),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf11b78b[1]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_a031887 (
    .a(al_6896ad14),
    .b(al_e4c850aa),
    .c(al_c289c50a[0]),
    .d(al_c289c50a[1]),
    .e(al_c289c50a[2]),
    .o(al_ce5f7b78));
  AL_DFF_0 al_64242e2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5699c1e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbeafa67[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    al_e1ac75ab (
    .a(al_10f0cebf),
    .b(al_cbeafa67[2]),
    .c(al_8ed48b41[2]),
    .d(al_18fc9355),
    .o(al_e5699c1e));
  AL_DFF_0 al_db0015d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_fd46e088[0]));
  AL_DFF_0 al_8ed8024f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_fd46e088[1]));
  AL_DFF_0 al_97b9705f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_d76fa964[2]));
  AL_DFF_0 al_689dab56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_57cd6e45[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_c289c50a[0]));
  AL_DFF_0 al_dbd8f608 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_57cd6e45[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_c289c50a[1]));
  AL_DFF_0 al_985e0e66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_57cd6e45[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_c289c50a[2]));
  AL_DFF_0 al_5d8c7dd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_90c83bf9[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_4a605a24[0]));
  AL_DFF_0 al_21e704d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_90c83bf9[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_4a605a24[1]));
  AL_DFF_0 al_7564e5bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_526d80ee[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b57d409[0]));
  AL_DFF_0 al_db811d4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_526d80ee[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b57d409[1]));
  AL_DFF_0 al_3e2d1382 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_526d80ee[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b57d409[2]));
  AL_DFF_0 al_3936e8d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_526d80ee[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b57d409[3]));
  AL_DFF_0 al_82948e72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_526d80ee[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b57d409[4]));
  AL_DFF_0 al_82fdea2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44b93047[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fc7c448b[0]));
  AL_DFF_0 al_8f693485 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44b93047[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fc7c448b[1]));
  AL_DFF_0 al_4ad94ea7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44b93047[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fc7c448b[2]));
  AL_DFF_0 al_b5ac5007 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44b93047[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fc7c448b[3]));
  AL_DFF_0 al_146dc4c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44b93047[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fc7c448b[4]));
  AL_DFF_0 al_dacb832d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f585ca5[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d206e68[0]));
  AL_DFF_0 al_8a9f25f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f585ca5[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d206e68[1]));
  AL_DFF_0 al_aef0c063 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f585ca5[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d206e68[2]));
  AL_DFF_0 al_6c8e8e8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f585ca5[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d206e68[3]));
  AL_DFF_0 al_5d62bc23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4f585ca5[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d206e68[4]));
  AL_DFF_0 al_20644e36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6ac4cff[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce0a0d6b[0]));
  AL_DFF_0 al_e70439b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6ac4cff[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce0a0d6b[1]));
  AL_DFF_0 al_7e505c33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6ac4cff[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce0a0d6b[2]));
  AL_DFF_0 al_c5879ae8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6ac4cff[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce0a0d6b[3]));
  AL_DFF_0 al_1cb96fb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6ac4cff[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce0a0d6b[4]));
  AL_DFF_0 al_ba4e19a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_afe3d62c[3]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_8278c32[3]));
  AL_DFF_0 al_1ed6f895 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_afe3d62c[4]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_8278c32[4]));
  AL_DFF_0 al_751b4d78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_afe3d62c[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_8278c32[0]));
  AL_DFF_0 al_7dd41a86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_afe3d62c[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_8278c32[1]));
  AL_DFF_0 al_51ca0d13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_afe3d62c[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_8278c32[2]));
  AL_DFF_0 al_2733f1f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[0]));
  AL_DFF_0 al_ee69f28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[1]));
  AL_DFF_0 al_ff347d22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[2]));
  AL_DFF_0 al_3bb4467f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[11]));
  AL_DFF_0 al_1f8d4526 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[12]));
  AL_DFF_0 al_98b95f7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[13]));
  AL_DFF_0 al_e53bf477 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[14]));
  AL_DFF_0 al_5e1e9b6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[15]));
  AL_DFF_0 al_292a3e31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[16]));
  AL_DFF_0 al_8daf454c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[17]));
  AL_DFF_0 al_3e3bce3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[24]));
  AL_DFF_0 al_562b47f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[25]));
  AL_DFF_0 al_2b7520e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[26]));
  AL_DFF_0 al_ffeb7e5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[27]));
  AL_DFF_0 al_5447371d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[28]));
  AL_DFF_0 al_cb6a4823 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[29]));
  AL_DFF_0 al_f7a8ddc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[30]));
  AL_DFF_0 al_90ab8947 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[31]));
  AL_DFF_0 al_5d0082ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[32]));
  AL_DFF_0 al_240b8546 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[33]));
  AL_DFF_0 al_b339da5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[34]));
  AL_DFF_0 al_e07b8600 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[35]));
  AL_DFF_0 al_b1411d8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[36]));
  AL_DFF_0 al_14c824af (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[37]));
  AL_DFF_0 al_7722fc87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[44]));
  AL_DFF_0 al_53c5d507 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[45]));
  AL_DFF_0 al_d95f80da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9af4975[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ed48b41[46]));
  AL_DFF_0 al_2af8687 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[0]));
  AL_DFF_0 al_25872e0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[1]));
  AL_DFF_0 al_378178b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[2]));
  AL_DFF_0 al_7fafef63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[11]));
  AL_DFF_0 al_e5dc2d5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[12]));
  AL_DFF_0 al_63a86ebc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[13]));
  AL_DFF_0 al_224aa500 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[14]));
  AL_DFF_0 al_711f56a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[15]));
  AL_DFF_0 al_1b2bd512 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[16]));
  AL_DFF_0 al_902efb92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[17]));
  AL_DFF_0 al_de1b61c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[24]));
  AL_DFF_0 al_be615abd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[25]));
  AL_DFF_0 al_bf0abe8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[26]));
  AL_DFF_0 al_ea853228 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[27]));
  AL_DFF_0 al_2122894c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[28]));
  AL_DFF_0 al_75a81ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[29]));
  AL_DFF_0 al_9b5c5ec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[30]));
  AL_DFF_0 al_f1543ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[31]));
  AL_DFF_0 al_e341b069 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[32]));
  AL_DFF_0 al_14ffb80e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[33]));
  AL_DFF_0 al_b1b04dbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[34]));
  AL_DFF_0 al_8f3b3115 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[35]));
  AL_DFF_0 al_b898f814 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[36]));
  AL_DFF_0 al_9be313eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[37]));
  AL_DFF_0 al_1f4c184f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[44]));
  AL_DFF_0 al_6cc8d10f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[45]));
  AL_DFF_0 al_3ab48cee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_f21eb389[0]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_1f1a358[46]));
  AL_DFF_0 al_f239c27f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[0]));
  AL_DFF_0 al_ca79ec47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[1]));
  AL_DFF_0 al_ddefe5a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[2]));
  AL_DFF_0 al_eab72e0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[11]));
  AL_DFF_0 al_a128d43c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[12]));
  AL_DFF_0 al_d608095f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[13]));
  AL_DFF_0 al_9f92ec33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[14]));
  AL_DFF_0 al_f4a5d4f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[15]));
  AL_DFF_0 al_b003e6c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[16]));
  AL_DFF_0 al_f086aca2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[17]));
  AL_DFF_0 al_de336d11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[24]));
  AL_DFF_0 al_11a29f59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[25]));
  AL_DFF_0 al_44ad53ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[26]));
  AL_DFF_0 al_1b2a37d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[27]));
  AL_DFF_0 al_f26b6181 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[28]));
  AL_DFF_0 al_ceadcd02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[29]));
  AL_DFF_0 al_5dbe6b9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[30]));
  AL_DFF_0 al_1cfe9d37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[31]));
  AL_DFF_0 al_2c849c5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[32]));
  AL_DFF_0 al_85f469d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[33]));
  AL_DFF_0 al_84afdd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[34]));
  AL_DFF_0 al_38418629 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[35]));
  AL_DFF_0 al_29c7123c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[36]));
  AL_DFF_0 al_9b9cde9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[37]));
  AL_DFF_0 al_ec6827f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[44]));
  AL_DFF_0 al_7587a89d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[45]));
  AL_DFF_0 al_cdac83c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_f21eb389[1]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_9840f3f[46]));
  AL_DFF_0 al_9958f5f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[0]));
  AL_DFF_0 al_d653936f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[1]));
  AL_DFF_0 al_677e8f0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[2]));
  AL_DFF_0 al_6964d8b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[11]));
  AL_DFF_0 al_84229964 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[12]));
  AL_DFF_0 al_4590b10b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[13]));
  AL_DFF_0 al_eb474d5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[14]));
  AL_DFF_0 al_3386d3d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[15]));
  AL_DFF_0 al_dc341f0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[16]));
  AL_DFF_0 al_cc6399ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[17]));
  AL_DFF_0 al_5b9d6cea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[24]));
  AL_DFF_0 al_940686d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[25]));
  AL_DFF_0 al_3e34c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[26]));
  AL_DFF_0 al_ba08dd9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[27]));
  AL_DFF_0 al_32dae184 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[28]));
  AL_DFF_0 al_c6764056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[29]));
  AL_DFF_0 al_6329aff3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[30]));
  AL_DFF_0 al_d60f6b74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[31]));
  AL_DFF_0 al_79916916 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[32]));
  AL_DFF_0 al_40af1be2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[33]));
  AL_DFF_0 al_1b5af3d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[34]));
  AL_DFF_0 al_5037ae03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[35]));
  AL_DFF_0 al_41f99be7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[36]));
  AL_DFF_0 al_2a2d3547 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[37]));
  AL_DFF_0 al_d8033bc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[44]));
  AL_DFF_0 al_724a68d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[45]));
  AL_DFF_0 al_ed0a5462 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_f21eb389[2]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7dc43980[46]));
  AL_DFF_0 al_4c40467c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[0]));
  AL_DFF_0 al_aed6973d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[1]));
  AL_DFF_0 al_20d0f43b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[2]));
  AL_DFF_0 al_f9d327e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[11]));
  AL_DFF_0 al_c35c84b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[12]));
  AL_DFF_0 al_d0243eb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[13]));
  AL_DFF_0 al_154c4de2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[14]));
  AL_DFF_0 al_8bd6c98d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[15]));
  AL_DFF_0 al_12212fa8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[16]));
  AL_DFF_0 al_789559f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[17]));
  AL_DFF_0 al_566c9702 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[24]));
  AL_DFF_0 al_6098e23b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[25]));
  AL_DFF_0 al_6dff732c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[26]));
  AL_DFF_0 al_71b73414 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[27]));
  AL_DFF_0 al_eb7ffa7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[28]));
  AL_DFF_0 al_e45d57d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[29]));
  AL_DFF_0 al_3beb38e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[30]));
  AL_DFF_0 al_c624f191 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[31]));
  AL_DFF_0 al_c1c0f7e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[32]));
  AL_DFF_0 al_2f1c6573 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[33]));
  AL_DFF_0 al_8c92ce34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[34]));
  AL_DFF_0 al_73c14532 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[35]));
  AL_DFF_0 al_c4ff3514 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[36]));
  AL_DFF_0 al_1e28f04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[37]));
  AL_DFF_0 al_531f00c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[44]));
  AL_DFF_0 al_fb34c9fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[45]));
  AL_DFF_0 al_55398e3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_f21eb389[3]),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_198cecf1[46]));
  AL_DFF_0 al_25c743a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bfcf9d28[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_bd042336[0]));
  AL_DFF_0 al_e5731491 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bfcf9d28[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_bd042336[1]));
  AL_DFF_0 al_8a38cdb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3612f044[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_66e5f5b5[0]));
  AL_DFF_0 al_939aebc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3612f044[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_66e5f5b5[1]));
  AL_DFF_0 al_53cc3b42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[0]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e42ac584[0]));
  AL_DFF_0 al_c16ff76e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[1]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e42ac584[1]));
  AL_DFF_0 al_bc995789 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[2]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e42ac584[2]));
  AL_DFF_0 al_b5eef862 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[3]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e42ac584[3]));
  AL_DFF_0 al_85d870ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[4]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e42ac584[4]));
  AL_DFF_0 al_19258cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[0]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_96dda245[0]));
  AL_DFF_0 al_99678e8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[1]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_96dda245[1]));
  AL_DFF_0 al_b6aa26dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[2]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_96dda245[2]));
  AL_DFF_0 al_21e73ac3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[3]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_96dda245[3]));
  AL_DFF_0 al_b19386e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[4]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_96dda245[4]));
  AL_DFF_0 al_25014e63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[0]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_535746d5[0]));
  AL_DFF_0 al_f1ec2ec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[1]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_535746d5[1]));
  AL_DFF_0 al_bc89f531 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[2]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_535746d5[2]));
  AL_DFF_0 al_75902a13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[3]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_535746d5[3]));
  AL_DFF_0 al_aaf2d9bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[4]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_535746d5[4]));
  AL_DFF_0 al_d1495a0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[0]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c8aa6814[0]));
  AL_DFF_0 al_240e448b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[1]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c8aa6814[1]));
  AL_DFF_0 al_67e98c99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[2]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c8aa6814[2]));
  AL_DFF_0 al_fcb19886 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[3]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c8aa6814[3]));
  AL_DFF_0 al_28110b85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8023991e[4]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c8aa6814[4]));
  AL_DFF_0 al_500f6071 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_14c34e2f[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_40b9c486[0]));
  AL_DFF_0 al_16e006a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_14c34e2f[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_40b9c486[1]));
  AL_DFF_0 al_c2abdd11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c8d0e932[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7a6f3e1[0]));
  AL_DFF_0 al_d0ff0df0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c8d0e932[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7a6f3e1[1]));
  AL_DFF_0 al_a30727ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c8d0e932[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7a6f3e1[2]));
  AL_DFF_0 al_301c6813 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c8d0e932[3]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_7a6f3e1[3]));
  AL_DFF_0 al_3c43296b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[0]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[0]));
  AL_DFF_0 al_e94ca64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[1]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[1]));
  AL_DFF_0 al_ed2f8f7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[2]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[2]));
  AL_DFF_0 al_8b548203 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[11]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[11]));
  AL_DFF_0 al_89b8d1f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[12]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[12]));
  AL_DFF_0 al_35128c40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[13]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[13]));
  AL_DFF_0 al_f328a994 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[14]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[14]));
  AL_DFF_0 al_9bbf47dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[15]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[15]));
  AL_DFF_0 al_95da2835 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[16]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[16]));
  AL_DFF_0 al_cc26dfd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[17]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[17]));
  AL_DFF_0 al_bca3a098 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[44]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[44]));
  AL_DFF_0 al_c34e7656 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[45]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[45]));
  AL_DFF_0 al_d27855ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[46]),
    .en(al_9119fd7[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8664dd36[46]));
  AL_DFF_0 al_f1810024 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[0]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[0]));
  AL_DFF_0 al_19bdbf90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[1]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[1]));
  AL_DFF_0 al_be56935d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[2]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[2]));
  AL_DFF_0 al_9ff121e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[11]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[11]));
  AL_DFF_0 al_fe5f41e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[12]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[12]));
  AL_DFF_0 al_f95db2fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[13]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[13]));
  AL_DFF_0 al_2933c00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[14]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[14]));
  AL_DFF_0 al_f685bffc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[15]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[15]));
  AL_DFF_0 al_5774b8f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[16]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[16]));
  AL_DFF_0 al_a0e007ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[17]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[17]));
  AL_DFF_0 al_1fe570a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[44]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[44]));
  AL_DFF_0 al_ba2a445e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[45]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[45]));
  AL_DFF_0 al_e569fd59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[46]),
    .en(al_9119fd7[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_393e4b3[46]));
  AL_DFF_0 al_e64d832 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[0]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[0]));
  AL_DFF_0 al_10682ee7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[1]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[1]));
  AL_DFF_0 al_8d9e0789 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[2]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[2]));
  AL_DFF_0 al_1d4f333d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[11]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[11]));
  AL_DFF_0 al_c7ccb85f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[12]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[12]));
  AL_DFF_0 al_d5803ae5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[13]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[13]));
  AL_DFF_0 al_7a9c0de8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[14]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[14]));
  AL_DFF_0 al_4e11ad80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[15]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[15]));
  AL_DFF_0 al_3f5f91c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[16]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[16]));
  AL_DFF_0 al_14d88bfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[17]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[17]));
  AL_DFF_0 al_6200b4f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[44]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[44]));
  AL_DFF_0 al_25990911 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[45]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[45]));
  AL_DFF_0 al_6c49a87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[46]),
    .en(al_9119fd7[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6ae1e35[46]));
  AL_DFF_0 al_4e76cd46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[0]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[0]));
  AL_DFF_0 al_ae3524ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[1]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[1]));
  AL_DFF_0 al_2a5951dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[2]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[2]));
  AL_DFF_0 al_f1c6128 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[11]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[11]));
  AL_DFF_0 al_d140169f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[12]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[12]));
  AL_DFF_0 al_e8fb3b69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[13]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[13]));
  AL_DFF_0 al_1733d03f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[14]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[14]));
  AL_DFF_0 al_b63782c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[15]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[15]));
  AL_DFF_0 al_27fe2ed9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[16]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[16]));
  AL_DFF_0 al_aa4802a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[17]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[17]));
  AL_DFF_0 al_9119c97e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[44]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[44]));
  AL_DFF_0 al_e523dc5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[45]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[45]));
  AL_DFF_0 al_fb9c5c16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8ed48b41[46]),
    .en(al_9119fd7[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b56343fc[46]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_ec04cd40 (
    .a(al_5b931dce),
    .b(al_fbe54a4d),
    .c(al_c289c50a[2]),
    .o(al_10f0cebf));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    al_502f042b (
    .a(al_10f0cebf),
    .b(al_8ed48b41[0]),
    .c(al_53bb123b[2]),
    .d(al_18fc9355),
    .o(al_e75d1e47));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    al_b1e3f702 (
    .a(al_10f0cebf),
    .b(al_8ed48b41[1]),
    .c(al_53bb123b[3]),
    .d(al_18fc9355),
    .o(al_7a20d1b6));
  AL_DFF_0 al_73db0e27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e75d1e47),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53bb123b[2]));
  AL_DFF_0 al_e0f641f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7a20d1b6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53bb123b[3]));
  AL_DFF_0 al_4d6d55c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b90e2b30[3]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_31a603ae[3]));
  AL_DFF_0 al_51a5cc7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b90e2b30[4]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_31a603ae[4]));
  AL_DFF_0 al_5bd6452f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b90e2b30[0]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_31a603ae[0]));
  AL_DFF_0 al_ec797870 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b90e2b30[1]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_31a603ae[1]));
  AL_DFF_0 al_cefd7ef5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b90e2b30[2]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_31a603ae[2]));
  AL_DFF_0 al_10b761d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[11]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2602b5cf[13]));
  AL_DFF_0 al_3c02c616 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[12]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2602b5cf[14]));
  AL_DFF_0 al_8a9cd5c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[13]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2602b5cf[15]));
  AL_DFF_0 al_8eff74fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[14]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2602b5cf[16]));
  AL_DFF_0 al_2cf0bd69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[15]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2602b5cf[17]));
  AL_DFF_0 al_f0a48654 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[16]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2602b5cf[18]));
  AL_DFF_0 al_53464fb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41f34c81[17]),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_2602b5cf[19]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b9fb6935 (
    .i(al_a3c26eaf),
    .o(al_2ccb9cac));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_332c4ffb (
    .i(al_2ccb9cac),
    .o(al_18fc9355));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*B*~(C)*D*E)"),
    .INIT(32'h0800fbcf))
    al_85b55c96 (
    .a(al_6e677e24),
    .b(al_c289c50a[0]),
    .c(al_c289c50a[1]),
    .d(al_c289c50a[2]),
    .e(al_8278c32[0]),
    .o(al_afe3d62c[0]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haacaa0aa))
    al_c48bfc46 (
    .a(al_637e5e2a[4]),
    .b(al_acf6f93e),
    .c(al_c289c50a[0]),
    .d(al_c289c50a[1]),
    .e(al_c289c50a[2]),
    .o(al_afe3d62c[4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_e6d4902a (
    .a(al_afe3d62c[4]),
    .b(al_afe3d62c[3]),
    .c(al_afe3d62c[2]),
    .d(al_afe3d62c[1]),
    .e(al_afe3d62c[0]),
    .o(al_69c0e2e6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~((F@E))+A*~(B)*~(C)*~(D)*~((F@E))+~(A)*B*~(C)*~(D)*~((F@E))+A*B*~(C)*~(D)*~((F@E))+~(A)*B*C*~(D)*~((F@E))+A*B*C*~(D)*~((F@E))+~(A)*~(B)*~(C)*D*~((F@E))+A*~(B)*~(C)*D*~((F@E))+A*B*~(C)*D*~((F@E))+~(A)*~(B)*C*D*~((F@E))+A*~(B)*C*D*~((F@E))+~(A)*B*C*D*~((F@E))+A*B*C*D*~((F@E))+A*B*~(C)*D*(F@E))"),
    .INIT(64'hfbcf08000800fbcf))
    al_1621631e (
    .a(al_d712b15f),
    .b(al_c289c50a[0]),
    .c(al_c289c50a[1]),
    .d(al_c289c50a[2]),
    .e(al_8278c32[0]),
    .f(al_8278c32[1]),
    .o(al_afe3d62c[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C@(~B*~A))"),
    .INIT(8'h1e))
    al_99035c0a (
    .a(al_8278c32[0]),
    .b(al_8278c32[1]),
    .c(al_8278c32[2]),
    .o(al_59c12bba));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55c55055))
    al_22981ea6 (
    .a(al_59c12bba),
    .b(al_fd39d17d),
    .c(al_c289c50a[0]),
    .d(al_c289c50a[1]),
    .e(al_c289c50a[2]),
    .o(al_afe3d62c[2]));
  AL_MAP_LUT4 #(
    .EQN("~(D@(~C*~B*~A))"),
    .INIT(16'h01fe))
    al_9507b958 (
    .a(al_8278c32[0]),
    .b(al_8278c32[1]),
    .c(al_8278c32[2]),
    .d(al_8278c32[3]),
    .o(al_19756cb7));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55c55055))
    al_4bd93db5 (
    .a(al_19756cb7),
    .b(al_112c6aa0),
    .c(al_c289c50a[0]),
    .d(al_c289c50a[1]),
    .e(al_c289c50a[2]),
    .o(al_afe3d62c[3]));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~C*~B*~A))"),
    .INIT(32'hfffe0001))
    al_2742bbbe (
    .a(al_8278c32[0]),
    .b(al_8278c32[1]),
    .c(al_8278c32[2]),
    .d(al_8278c32[3]),
    .e(al_8278c32[4]),
    .o(al_637e5e2a[4]));
  AL_DFF_0 al_978bc18f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69c0e2e6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ca5b8a7));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_f4ce1f61 (
    .a(al_58d81d6c),
    .b(al_66e5f5b5[0]),
    .o(al_3612f044[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    al_78c1e047 (
    .a(al_58d81d6c),
    .b(al_66e5f5b5[0]),
    .c(al_66e5f5b5[1]),
    .o(al_3612f044[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_b5e791fc (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_3612f044[0]),
    .d(al_3612f044[1]),
    .o(al_15aa8dca));
  AL_DFF_0 al_506a0d33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_15aa8dca),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_23659fe5));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_7b202978 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[5]),
    .c(al_1f1a358[0]),
    .o(al_cabc97d1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a2ebbd89 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[5]),
    .c(al_9840f3f[0]),
    .o(al_16a767cd[0]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1893c360 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[5]),
    .c(al_7dc43980[0]),
    .o(al_42da1f0d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4c1d5ad1 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[5]),
    .c(al_198cecf1[0]),
    .o(al_17da2162[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_74477219 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_cabc97d1),
    .d(al_42da1f0d),
    .e(al_16a767cd[0]),
    .f(al_17da2162[0]),
    .o(al_d9af4975[0]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_fd397566 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[6]),
    .c(al_1f1a358[11]),
    .o(al_4a355d24));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e0fa2110 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[6]),
    .c(al_9840f3f[11]),
    .o(al_16a767cd[11]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_2bcaaeca (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[6]),
    .c(al_7dc43980[11]),
    .o(al_12d74399));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_23daf7da (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[6]),
    .c(al_198cecf1[11]),
    .o(al_17da2162[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_2bf02fe7 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_4a355d24),
    .d(al_12d74399),
    .e(al_16a767cd[11]),
    .f(al_17da2162[11]),
    .o(al_d9af4975[11]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_48a9db05 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[7]),
    .c(al_1f1a358[12]),
    .o(al_ce2d52c6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e2c6b7f (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[7]),
    .c(al_9840f3f[12]),
    .o(al_16a767cd[12]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_3f090dfd (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[7]),
    .c(al_7dc43980[12]),
    .o(al_c3834b72));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2040bb7 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[7]),
    .c(al_198cecf1[12]),
    .o(al_17da2162[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_7ac9bcd5 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_ce2d52c6),
    .d(al_c3834b72),
    .e(al_16a767cd[12]),
    .f(al_17da2162[12]),
    .o(al_d9af4975[12]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f4277f81 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[8]),
    .c(al_1f1a358[13]),
    .o(al_ac6ac5f3));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e71dd2a4 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[8]),
    .c(al_9840f3f[13]),
    .o(al_16a767cd[13]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e864493f (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[8]),
    .c(al_7dc43980[13]),
    .o(al_553348a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_81e83856 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[8]),
    .c(al_198cecf1[13]),
    .o(al_17da2162[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_bab86f0e (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_ac6ac5f3),
    .d(al_553348a),
    .e(al_16a767cd[13]),
    .f(al_17da2162[13]),
    .o(al_d9af4975[13]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b88de295 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[9]),
    .c(al_7dc43980[14]),
    .o(al_709c747d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_362a7808 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[9]),
    .c(al_198cecf1[14]),
    .o(al_17da2162[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_788f868a (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[9]),
    .c(al_9840f3f[14]),
    .o(al_16a767cd[14]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_5f6de536 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[9]),
    .c(al_1f1a358[14]),
    .o(al_c7d91c95));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haebf26378c9d0415))
    al_2eb83b4c (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_709c747d),
    .d(al_c7d91c95),
    .e(al_17da2162[14]),
    .f(al_16a767cd[14]),
    .o(al_d9af4975[14]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a53e0fd2 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[10]),
    .c(al_1f1a358[15]),
    .o(al_a27e626a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e6e1885c (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[10]),
    .c(al_9840f3f[15]),
    .o(al_16a767cd[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_173c357c (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[10]),
    .c(al_7dc43980[15]),
    .o(al_9bbc19f6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_df5ea44a (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[10]),
    .c(al_198cecf1[15]),
    .o(al_17da2162[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_dadcedc6 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_a27e626a),
    .d(al_9bbc19f6),
    .e(al_16a767cd[15]),
    .f(al_17da2162[15]),
    .o(al_d9af4975[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_bf5f1d1f (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[11]),
    .c(al_1f1a358[16]),
    .o(al_3e8e72a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_84d8dcc0 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[11]),
    .c(al_9840f3f[16]),
    .o(al_16a767cd[16]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d51d9473 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[11]),
    .c(al_7dc43980[16]),
    .o(al_8c4b2a57));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d039f86b (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[11]),
    .c(al_198cecf1[16]),
    .o(al_17da2162[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_940c6c09 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_3e8e72a),
    .d(al_8c4b2a57),
    .e(al_16a767cd[16]),
    .f(al_17da2162[16]),
    .o(al_d9af4975[16]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_cbae0e4b (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[12]),
    .c(al_1f1a358[17]),
    .o(al_6e29173f));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4f7efb58 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[12]),
    .c(al_9840f3f[17]),
    .o(al_16a767cd[17]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d33165dd (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[12]),
    .c(al_7dc43980[17]),
    .o(al_ce965e5b));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f21ff470 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[12]),
    .c(al_198cecf1[17]),
    .o(al_17da2162[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_ba6d8ddd (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_6e29173f),
    .d(al_ce965e5b),
    .e(al_16a767cd[17]),
    .f(al_17da2162[17]),
    .o(al_d9af4975[17]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d1d4ab2b (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[3]),
    .c(al_1f1a358[1]),
    .o(al_1cc0dee2));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d2f12c96 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[3]),
    .c(al_9840f3f[1]),
    .o(al_16a767cd[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_46dd4aba (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[3]),
    .c(al_7dc43980[1]),
    .o(al_e2e9d990));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8791c943 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[3]),
    .c(al_198cecf1[1]),
    .o(al_17da2162[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_a8ba93ea (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_1cc0dee2),
    .d(al_e2e9d990),
    .e(al_16a767cd[1]),
    .f(al_17da2162[1]),
    .o(al_d9af4975[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_7059a7d8 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[13]),
    .c(al_1f1a358[24]),
    .o(al_c56838c1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_72878894 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[13]),
    .c(al_9840f3f[24]),
    .o(al_16a767cd[24]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_93db4db6 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[13]),
    .c(al_7dc43980[24]),
    .o(al_5abac53e));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1d77381c (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[13]),
    .c(al_198cecf1[24]),
    .o(al_17da2162[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_603a6e0f (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_c56838c1),
    .d(al_5abac53e),
    .e(al_16a767cd[24]),
    .f(al_17da2162[24]),
    .o(al_d9af4975[24]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1f11c9de (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[14]),
    .c(al_1f1a358[25]),
    .o(al_a89a7f53));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8fde3893 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[14]),
    .c(al_9840f3f[25]),
    .o(al_16a767cd[25]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_41a0b255 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[14]),
    .c(al_7dc43980[25]),
    .o(al_d62c6586));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_57805a44 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[14]),
    .c(al_198cecf1[25]),
    .o(al_17da2162[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_93a3de48 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_a89a7f53),
    .d(al_d62c6586),
    .e(al_16a767cd[25]),
    .f(al_17da2162[25]),
    .o(al_d9af4975[25]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f8777232 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[15]),
    .c(al_1f1a358[26]),
    .o(al_4b666b4a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fa31aa0f (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[15]),
    .c(al_9840f3f[26]),
    .o(al_16a767cd[26]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_682b8a81 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[15]),
    .c(al_7dc43980[26]),
    .o(al_ac02de78));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4b9c961f (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[15]),
    .c(al_198cecf1[26]),
    .o(al_17da2162[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_6a7cb6f7 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_4b666b4a),
    .d(al_ac02de78),
    .e(al_16a767cd[26]),
    .f(al_17da2162[26]),
    .o(al_d9af4975[26]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_365409d2 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[16]),
    .c(al_1f1a358[27]),
    .o(al_ba842b48));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f9a72447 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[16]),
    .c(al_9840f3f[27]),
    .o(al_16a767cd[27]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b14f510e (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[16]),
    .c(al_7dc43980[27]),
    .o(al_aefc71a0));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bd861f2c (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[16]),
    .c(al_198cecf1[27]),
    .o(al_17da2162[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_4b1fcad4 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_ba842b48),
    .d(al_aefc71a0),
    .e(al_16a767cd[27]),
    .f(al_17da2162[27]),
    .o(al_d9af4975[27]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_4763ab6b (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[17]),
    .c(al_1f1a358[28]),
    .o(al_5feeb4d9));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_924f8ca0 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[17]),
    .c(al_9840f3f[28]),
    .o(al_16a767cd[28]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b200c456 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[17]),
    .c(al_7dc43980[28]),
    .o(al_4b633b4a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_652788ab (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[17]),
    .c(al_198cecf1[28]),
    .o(al_17da2162[28]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_287589f6 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_5feeb4d9),
    .d(al_4b633b4a),
    .e(al_16a767cd[28]),
    .f(al_17da2162[28]),
    .o(al_d9af4975[28]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d2bf64d0 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[18]),
    .c(al_1f1a358[29]),
    .o(al_db625dc2));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_26a700b3 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[18]),
    .c(al_9840f3f[29]),
    .o(al_16a767cd[29]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_64eb12c2 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[18]),
    .c(al_7dc43980[29]),
    .o(al_f15041ee));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ad4f9638 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[18]),
    .c(al_198cecf1[29]),
    .o(al_17da2162[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_fd964232 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_db625dc2),
    .d(al_f15041ee),
    .e(al_16a767cd[29]),
    .f(al_17da2162[29]),
    .o(al_d9af4975[29]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a13020ed (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[4]),
    .c(al_1f1a358[2]),
    .o(al_42951d78));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5a1c907c (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[4]),
    .c(al_9840f3f[2]),
    .o(al_16a767cd[2]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e35d8f25 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[4]),
    .c(al_7dc43980[2]),
    .o(al_1ca1a962));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b2743d90 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[4]),
    .c(al_198cecf1[2]),
    .o(al_17da2162[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_841c96e8 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_42951d78),
    .d(al_1ca1a962),
    .e(al_16a767cd[2]),
    .f(al_17da2162[2]),
    .o(al_d9af4975[2]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_8eba6b63 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[19]),
    .c(al_1f1a358[30]),
    .o(al_b3e959dd));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fe49c6d5 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[19]),
    .c(al_9840f3f[30]),
    .o(al_16a767cd[30]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e5aaf7ab (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[19]),
    .c(al_7dc43980[30]),
    .o(al_b7cccbae));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5678c0dd (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[19]),
    .c(al_198cecf1[30]),
    .o(al_17da2162[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_9c0b4b71 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_b3e959dd),
    .d(al_b7cccbae),
    .e(al_16a767cd[30]),
    .f(al_17da2162[30]),
    .o(al_d9af4975[30]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_afb6d238 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[20]),
    .c(al_1f1a358[31]),
    .o(al_d6b1e9ef));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ce3b7fd2 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[20]),
    .c(al_9840f3f[31]),
    .o(al_16a767cd[31]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_4831953d (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[20]),
    .c(al_7dc43980[31]),
    .o(al_cff520de));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c976d201 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[20]),
    .c(al_198cecf1[31]),
    .o(al_17da2162[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_31188236 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_d6b1e9ef),
    .d(al_cff520de),
    .e(al_16a767cd[31]),
    .f(al_17da2162[31]),
    .o(al_d9af4975[31]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_92eebb4d (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[21]),
    .c(al_1f1a358[32]),
    .o(al_709efed6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5782d426 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[21]),
    .c(al_9840f3f[32]),
    .o(al_16a767cd[32]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_fd248630 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[21]),
    .c(al_7dc43980[32]),
    .o(al_41779a5c));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ae731eee (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[21]),
    .c(al_198cecf1[32]),
    .o(al_17da2162[32]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_9c27f10f (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_709efed6),
    .d(al_41779a5c),
    .e(al_16a767cd[32]),
    .f(al_17da2162[32]),
    .o(al_d9af4975[32]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_80c82047 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[22]),
    .c(al_1f1a358[33]),
    .o(al_ec69184c));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3695634f (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[22]),
    .c(al_9840f3f[33]),
    .o(al_16a767cd[33]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6281f22f (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[22]),
    .c(al_7dc43980[33]),
    .o(al_bba532bd));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4e95a6f (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[22]),
    .c(al_198cecf1[33]),
    .o(al_17da2162[33]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_9adf2939 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_ec69184c),
    .d(al_bba532bd),
    .e(al_16a767cd[33]),
    .f(al_17da2162[33]),
    .o(al_d9af4975[33]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_7f1c8fad (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[23]),
    .c(al_1f1a358[34]),
    .o(al_12c68610));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_88a2a662 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[23]),
    .c(al_9840f3f[34]),
    .o(al_16a767cd[34]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d5e9abfd (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[23]),
    .c(al_7dc43980[34]),
    .o(al_59d2fcf));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_887f2881 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[23]),
    .c(al_198cecf1[34]),
    .o(al_17da2162[34]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_4f401f04 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_12c68610),
    .d(al_59d2fcf),
    .e(al_16a767cd[34]),
    .f(al_17da2162[34]),
    .o(al_d9af4975[34]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6e87d12b (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[24]),
    .c(al_1f1a358[35]),
    .o(al_7ff14cde));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_43f5a05f (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[24]),
    .c(al_9840f3f[35]),
    .o(al_16a767cd[35]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f74f9451 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[24]),
    .c(al_7dc43980[35]),
    .o(al_9b7ed9ba));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_69a9450e (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[24]),
    .c(al_198cecf1[35]),
    .o(al_17da2162[35]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_5f8409dc (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_7ff14cde),
    .d(al_9b7ed9ba),
    .e(al_16a767cd[35]),
    .f(al_17da2162[35]),
    .o(al_d9af4975[35]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6e95ba03 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[25]),
    .c(al_1f1a358[36]),
    .o(al_324d8fba));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ee2b16cc (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[25]),
    .c(al_9840f3f[36]),
    .o(al_16a767cd[36]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_37376a7f (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[25]),
    .c(al_7dc43980[36]),
    .o(al_af37d5e4));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3d4e1d1d (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[25]),
    .c(al_198cecf1[36]),
    .o(al_17da2162[36]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_b3390209 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_324d8fba),
    .d(al_af37d5e4),
    .e(al_16a767cd[36]),
    .f(al_17da2162[36]),
    .o(al_d9af4975[36]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_adb520e8 (
    .a(al_f21eb389[0]),
    .b(al_58fb4752[26]),
    .c(al_1f1a358[37]),
    .o(al_3799028a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5fa4b0b8 (
    .a(al_f21eb389[1]),
    .b(al_58fb4752[26]),
    .c(al_9840f3f[37]),
    .o(al_16a767cd[37]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6f6e74f5 (
    .a(al_f21eb389[2]),
    .b(al_58fb4752[26]),
    .c(al_7dc43980[37]),
    .o(al_72d179c3));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4e4d751 (
    .a(al_f21eb389[3]),
    .b(al_58fb4752[26]),
    .c(al_198cecf1[37]),
    .o(al_17da2162[37]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_6ef70d3f (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_3799028a),
    .d(al_72d179c3),
    .e(al_16a767cd[37]),
    .f(al_17da2162[37]),
    .o(al_d9af4975[37]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_540b0fd0 (
    .a(al_f21eb389[0]),
    .b(al_88a8db2c[0]),
    .c(al_1f1a358[44]),
    .o(al_bb5bd57a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6247cbd9 (
    .a(al_f21eb389[1]),
    .b(al_88a8db2c[0]),
    .c(al_9840f3f[44]),
    .o(al_16a767cd[44]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6c8a6ce (
    .a(al_f21eb389[2]),
    .b(al_88a8db2c[0]),
    .c(al_7dc43980[44]),
    .o(al_9e317c87));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e5acf7b5 (
    .a(al_f21eb389[3]),
    .b(al_88a8db2c[0]),
    .c(al_198cecf1[44]),
    .o(al_17da2162[44]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_a9eb81a2 (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_bb5bd57a),
    .d(al_9e317c87),
    .e(al_16a767cd[44]),
    .f(al_17da2162[44]),
    .o(al_d9af4975[44]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_cd60ea56 (
    .a(al_f21eb389[0]),
    .b(al_88a8db2c[1]),
    .c(al_1f1a358[45]),
    .o(al_fd9fbb70));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2c92b321 (
    .a(al_f21eb389[1]),
    .b(al_88a8db2c[1]),
    .c(al_9840f3f[45]),
    .o(al_16a767cd[45]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_96a26fba (
    .a(al_f21eb389[2]),
    .b(al_88a8db2c[1]),
    .c(al_7dc43980[45]),
    .o(al_978813a6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6a51c4ce (
    .a(al_f21eb389[3]),
    .b(al_88a8db2c[1]),
    .c(al_198cecf1[45]),
    .o(al_17da2162[45]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_91c6362a (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_fd9fbb70),
    .d(al_978813a6),
    .e(al_16a767cd[45]),
    .f(al_17da2162[45]),
    .o(al_d9af4975[45]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7491b26c (
    .a(al_3612f044[0]),
    .b(al_66e5f5b5[1]),
    .o(al_f21eb389[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_424956e5 (
    .a(al_f21eb389[3]),
    .b(al_88a8db2c[2]),
    .c(al_198cecf1[46]),
    .o(al_17da2162[46]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_964c8c3e (
    .a(al_bfcf9d28[0]),
    .b(al_bfcf9d28[1]),
    .c(al_4f79a2d4),
    .d(al_9ea1824f),
    .e(al_16a767cd[46]),
    .f(al_17da2162[46]),
    .o(al_d9af4975[46]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_1c420802 (
    .a(al_3612f044[0]),
    .b(al_3612f044[1]),
    .o(al_f21eb389[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_d2decc00 (
    .a(al_3612f044[0]),
    .b(al_3612f044[1]),
    .o(al_f21eb389[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_7cae20eb (
    .a(al_3612f044[0]),
    .b(al_66e5f5b5[1]),
    .o(al_f21eb389[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ad79cc1 (
    .a(al_f21eb389[0]),
    .b(al_88a8db2c[2]),
    .c(al_1f1a358[46]),
    .o(al_4f79a2d4));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_549fbce0 (
    .a(al_f21eb389[1]),
    .b(al_88a8db2c[2]),
    .c(al_9840f3f[46]),
    .o(al_16a767cd[46]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_2b44d35f (
    .a(al_f21eb389[2]),
    .b(al_88a8db2c[2]),
    .c(al_7dc43980[46]),
    .o(al_9ea1824f));
  AL_DFF_0 al_7d836dfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2182cd10),
    .en(1'b1),
    .sr(al_18fc9355),
    .ss(1'b0),
    .q(al_891497d5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_50fabf2 (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[0]),
    .d(al_393e4b3[0]),
    .e(al_c6ae1e35[0]),
    .f(al_b56343fc[0]),
    .o(al_61973ebe));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_b20a7f5a (
    .a(al_c289c50a[0]),
    .b(al_c289c50a[1]),
    .o(al_fbe54a4d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_f8556c95 (
    .a(al_46fc25e7),
    .b(al_fb20038d),
    .c(al_1f586c30),
    .d(al_4ce39135),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_66395a07));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_62599ede (
    .a(al_627e01b),
    .b(al_58f4bcca),
    .c(al_a5fb3197),
    .d(al_865e3224),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_a23768c8));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_195601f0 (
    .a(al_fe185597),
    .b(al_f0cf2c1b),
    .c(al_b797198c),
    .d(al_8b71d8b7),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_be15f9bd));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_b2adf055 (
    .a(al_1ea50fd5),
    .b(al_48347124),
    .c(al_67f78c15),
    .d(al_3b14a515),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_646e2f99));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_abb550aa (
    .a(al_af3a3adf),
    .b(al_9384d2a6),
    .c(al_5c212f53),
    .d(al_d8c260df),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_d2a4a6b0));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_1cef336c (
    .a(al_cf63226f),
    .b(al_a0f44394),
    .c(al_73f87281),
    .d(al_79ca7989),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_82bab79d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_e2802b2 (
    .a(al_22d551b1),
    .b(al_ffaa6ed4),
    .c(al_f53cd64f),
    .d(al_b93ffb04),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_17c7de95));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_4c43d754 (
    .a(al_88d2570b),
    .b(al_ae9de7f7),
    .c(al_8ed48b41[0]),
    .o(al_45251641));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_d9c66a0d (
    .a(al_45251641),
    .b(al_cafe0ec3),
    .c(al_3c683e0a),
    .d(al_8ed48b41[0]),
    .e(al_8ed48b41[1]),
    .f(al_8ed48b41[31]),
    .o(al_11b8e521));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_103d8bc1 (
    .a(al_80336d41),
    .b(al_5bb79c4f),
    .c(al_b6b9db4),
    .d(al_42cfbe9b),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_3b042d56));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_901ce7ab (
    .a(al_61973ebe),
    .b(al_e4c850aa),
    .c(al_8ed48b41[0]),
    .o(al_41f34c81[0]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_5a25e07c (
    .a(al_cf05798c),
    .b(al_ddc7a73f),
    .c(al_8ed48b41[0]),
    .o(al_514e3a7));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_e7791fd7 (
    .a(al_514e3a7),
    .b(al_a620188b),
    .c(al_79ced939),
    .d(al_8ed48b41[0]),
    .e(al_8ed48b41[1]),
    .f(al_8ed48b41[33]),
    .o(al_ff98656b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_bfdbc1cb (
    .a(al_868dabaf),
    .b(al_25fc271e),
    .c(al_81d476eb),
    .d(al_699f3bb8),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_ef7c15ad));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_14d2890b (
    .a(al_7aadf07),
    .b(al_b7e2e71f),
    .c(al_8ed48b41[0]),
    .o(al_786b0491));
  AL_MAP_LUT6 #(
    .EQN("(F@~(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'hf0cc55550f33aaaa))
    al_b023495a (
    .a(al_786b0491),
    .b(al_5cd3a57d),
    .c(al_b2200d60),
    .d(al_8ed48b41[0]),
    .e(al_8ed48b41[1]),
    .f(al_8ed48b41[36]),
    .o(al_5a2ac1a2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_acff8de2 (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[1]),
    .d(al_393e4b3[1]),
    .e(al_c6ae1e35[1]),
    .f(al_b56343fc[1]),
    .o(al_f8db84b7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_34670610 (
    .a(al_ab1b96f9),
    .b(al_c34f057a),
    .c(al_fccfd8ff),
    .d(al_be66ece6),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_d77bb542));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_3e8c2416 (
    .a(al_9a04ce8f),
    .b(al_4c783ffb),
    .c(al_8ed48b41[0]),
    .o(al_9dfaf151));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_7e8cfae6 (
    .a(al_9dfaf151),
    .b(al_38c33a99),
    .c(al_310a635),
    .d(al_8ed48b41[0]),
    .e(al_8ed48b41[1]),
    .f(al_8ed48b41[35]),
    .o(al_c621ceb7));
  AL_MAP_LUT6 #(
    .EQN("((F@C)*(E@B)*(D@A))"),
    .INIT(64'h0102040810204080))
    al_a59e95e9 (
    .a(al_66395a07),
    .b(al_17c7de95),
    .c(al_3b042d56),
    .d(al_8ed48b41[25]),
    .e(al_8ed48b41[26]),
    .f(al_8ed48b41[28]),
    .o(al_6f281a7f));
  AL_MAP_LUT6 #(
    .EQN("(~B*A*(E@D)*(F@C))"),
    .INIT(64'h0002020000202000))
    al_baaf7e9a (
    .a(al_5a2ac1a2),
    .b(al_c621ceb7),
    .c(al_646e2f99),
    .d(al_82bab79d),
    .e(al_8ed48b41[30]),
    .f(al_8ed48b41[32]),
    .o(al_8d6dd847));
  AL_MAP_LUT6 #(
    .EQN("((D@C)*(E@B)*(F@A))"),
    .INIT(64'h0110044002200880))
    al_b7000174 (
    .a(al_be15f9bd),
    .b(al_d2a4a6b0),
    .c(al_ef7c15ad),
    .d(al_8ed48b41[24]),
    .e(al_8ed48b41[27]),
    .f(al_8ed48b41[29]),
    .o(al_d94dff22));
  AL_MAP_LUT6 #(
    .EQN("(~B*~A*(F@D)*(E@C))"),
    .INIT(64'h0001001001001000))
    al_e887e45e (
    .a(al_11b8e521),
    .b(al_ff98656b),
    .c(al_a23768c8),
    .d(al_d77bb542),
    .e(al_8ed48b41[34]),
    .f(al_8ed48b41[37]),
    .o(al_f22292ec));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_7d9288a6 (
    .a(al_b56598d),
    .b(al_122466dd),
    .c(al_195fd12),
    .d(al_91e55879),
    .e(al_8ed48b41[0]),
    .f(al_8ed48b41[1]),
    .o(al_4db2fe90));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*~B))"),
    .INIT(16'h0405))
    al_ff74fa30 (
    .a(al_4db2fe90),
    .b(al_58d81d6c),
    .c(al_25e1cc7),
    .d(al_23659fe5),
    .o(al_ef2f822e));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_535e7b77 (
    .a(al_8d6dd847),
    .b(al_f22292ec),
    .c(al_6f281a7f),
    .d(al_d94dff22),
    .e(al_ef2f822e),
    .f(al_fbe54a4d),
    .o(al_75fd0159));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(E*C*B*~A))"),
    .INIT(32'h00bf00ff))
    al_d950ddd8 (
    .a(al_25e1cc7),
    .b(al_c289c50a[0]),
    .c(al_c289c50a[1]),
    .d(al_c289c50a[2]),
    .e(al_c360bf4c[1]),
    .o(al_437081f2));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_b1e7cecf (
    .a(al_f8db84b7),
    .b(al_e4c850aa),
    .c(al_8ed48b41[1]),
    .o(al_41f34c81[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_88a1cda9 (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[45]),
    .d(al_393e4b3[45]),
    .e(al_c6ae1e35[45]),
    .f(al_b56343fc[45]),
    .o(al_f6e750ed));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_fe3dfd60 (
    .a(al_f6e750ed),
    .b(al_e4c850aa),
    .c(al_8ed48b41[45]),
    .o(al_f735a538));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_64414c8b (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[46]),
    .d(al_393e4b3[46]),
    .e(al_c6ae1e35[46]),
    .f(al_b56343fc[46]),
    .o(al_bf156068));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_be3a6e4e (
    .a(al_bf156068),
    .b(al_e4c850aa),
    .c(al_8ed48b41[46]),
    .o(al_41f34c81[46]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_2892d355 (
    .a(al_40b9c486[0]),
    .b(al_40b9c486[1]),
    .c(al_8664dd36[44]),
    .d(al_393e4b3[44]),
    .e(al_c6ae1e35[44]),
    .f(al_b56343fc[44]),
    .o(al_6158c618));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_41138ac6 (
    .a(al_6158c618),
    .b(al_e4c850aa),
    .c(al_8ed48b41[44]),
    .o(al_c9ddcee1));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_f85f05ac (
    .a(init_calib_complete),
    .b(al_90d84dc7[1]),
    .c(al_61f44420),
    .d(ddr_app_rdy),
    .o(al_58d81d6c));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d48ad5e7 (
    .a(al_41f34c81[46]),
    .b(al_c9ddcee1),
    .o(al_cd0bc85d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_29382551 (
    .a(al_41f34c81[0]),
    .b(al_41f34c81[1]),
    .c(al_51ceabf0),
    .d(al_3fdd9bd4),
    .e(al_724e96cb),
    .f(al_f6cbc027),
    .o(al_7b63babf));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~(~D*~(C*~A))))"),
    .INIT(32'h00233333))
    al_74f4e9f9 (
    .a(al_75fd0159),
    .b(al_7b63babf),
    .c(al_437081f2),
    .d(al_786dc891),
    .e(al_e4c850aa),
    .o(al_c20a9a7e));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_36a33bd (
    .a(al_cd0bc85d),
    .b(al_f735a538),
    .o(al_56be2a2c));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_7cf803b0 (
    .a(al_f735a538),
    .b(al_41f34c81[46]),
    .c(al_c9ddcee1),
    .d(al_4a605a24[0]),
    .e(al_4a605a24[1]),
    .o(al_f66d7bc0));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~(C*~B*A)))"),
    .INIT(32'h00ff0020))
    al_a26f4e6d (
    .a(al_c20a9a7e),
    .b(al_56be2a2c),
    .c(al_f66d7bc0),
    .d(al_b4c6b3bd),
    .e(al_891497d5),
    .o(al_2182cd10));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    al_a756f3c8 (
    .a(al_25e1cc7),
    .b(al_c289c50a[0]),
    .c(al_c289c50a[1]),
    .d(al_c289c50a[2]),
    .o(al_786dc891));
  AL_DFF_0 al_8f67709b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_40276cd4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90d84dc7[2]));
  AL_DFF_0 al_5f107ce5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8d431b3f),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_15ca36a));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_300df508 (
    .a(al_9860067e),
    .b(al_ad9637b9),
    .o(al_a0789cd8));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(~D*(A*C*~(E)*~(F)+A*C*~(E)*F+~(A)*~(C)*E*F+A*~(C)*E*F)))"),
    .INIT(64'h3330331333333313))
    al_34734637 (
    .a(al_114b0fe8),
    .b(al_15ca36a),
    .c(al_369e229d[0]),
    .d(al_369e229d[1]),
    .e(al_369e229d[2]),
    .f(al_f7e9a10b),
    .o(al_630da3b0));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_c4a4d8ec (
    .a(al_630da3b0),
    .b(al_c360bf4c[2]),
    .o(al_8d431b3f));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_d67c51d8 (
    .a(al_8941a5fb[0]),
    .b(al_8941a5fb[1]),
    .c(al_413c0926[0]),
    .d(al_59b0cd05[0]),
    .e(al_59b0cd05[1]),
    .o(al_cfa51fb3[0]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_a9c4fc30 (
    .a(al_8941a5fb[0]),
    .b(al_8941a5fb[1]),
    .c(al_413c0926[3]),
    .d(al_51cc7f19[0]),
    .e(al_51cc7f19[1]),
    .o(al_cfa51fb3[3]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_5cb37d54 (
    .a(al_8941a5fb[0]),
    .b(al_8941a5fb[1]),
    .c(al_413c0926[1]),
    .d(al_e9ebbe15[0]),
    .e(al_e9ebbe15[1]),
    .o(al_cfa51fb3[1]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(D*~(F@C)*~(E@B)))"),
    .INIT(64'h1555455551555455))
    al_9c408748 (
    .a(al_cfa51fb3[3]),
    .b(al_8941a5fb[0]),
    .c(al_8941a5fb[1]),
    .d(al_413c0926[2]),
    .e(al_c5c971b[0]),
    .f(al_c5c971b[1]),
    .o(al_94f083a0));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_c8ca174c (
    .a(al_94f083a0),
    .b(al_cfa51fb3[0]),
    .c(al_cfa51fb3[1]),
    .o(al_ca418906));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_f5694d02 (
    .a(al_ca418906),
    .b(al_a0789cd8),
    .c(al_c711503f),
    .o(al_114b0fe8));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*~A))"),
    .INIT(8'hc9))
    al_6ed2b368 (
    .a(al_1d36bc6d),
    .b(al_b0fb8887),
    .c(al_19e106e3),
    .o(al_21bd4e5d[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(~D*~B*~A))"),
    .INIT(16'hf0e1))
    al_eefd279b (
    .a(al_1d36bc6d),
    .b(al_b0fb8887),
    .c(al_a9552c76),
    .d(al_19e106e3),
    .o(al_21bd4e5d[2]));
  AL_MAP_LUT6 #(
    .EQN("(E@(~F*~D*~C*~B*~A))"),
    .INIT(64'hffff0000fffe0001))
    al_bc84fd8c (
    .a(al_1d36bc6d),
    .b(al_b0fb8887),
    .c(al_a9552c76),
    .d(al_4331638),
    .e(al_2a6634d6),
    .f(al_19e106e3),
    .o(al_21bd4e5d[4]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_d91e93ce (
    .a(al_1d36bc6d),
    .b(al_19e106e3),
    .o(al_21bd4e5d[0]));
  AL_MAP_LUT5 #(
    .EQN("(D@(~E*~C*~B*~A))"),
    .INIT(32'hff00fe01))
    al_4830f602 (
    .a(al_1d36bc6d),
    .b(al_b0fb8887),
    .c(al_a9552c76),
    .d(al_4331638),
    .e(al_19e106e3),
    .o(al_21bd4e5d[3]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_d0faf796 (
    .a(al_21bd4e5d[3]),
    .b(al_21bd4e5d[0]),
    .c(al_b0fb8887),
    .d(al_a9552c76),
    .e(al_2a6634d6),
    .o(al_61614b33[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_d9e78513 (
    .a(al_61614b33[0]),
    .b(al_19e106e3),
    .o(al_4bc24ece[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_32f09359 (
    .a(al_ac18355b[0]),
    .b(al_d0a384c4[0]),
    .c(al_1e043bfe[0]),
    .d(al_b0a8403e[0]),
    .e(al_11a7c870[0]),
    .f(al_11a7c870[1]),
    .o(al_3e345b21[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_eda06ffc (
    .a(al_ac18355b[1]),
    .b(al_d0a384c4[1]),
    .c(al_1e043bfe[1]),
    .d(al_b0a8403e[1]),
    .e(al_11a7c870[0]),
    .f(al_11a7c870[1]),
    .o(al_3e345b21[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_4fdfe072 (
    .a(al_ac18355b[2]),
    .b(al_d0a384c4[2]),
    .c(al_1e043bfe[2]),
    .d(al_b0a8403e[2]),
    .e(al_11a7c870[0]),
    .f(al_11a7c870[1]),
    .o(al_3e345b21[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_c41228f3 (
    .a(al_ac18355b[3]),
    .b(al_d0a384c4[3]),
    .c(al_1e043bfe[3]),
    .d(al_b0a8403e[3]),
    .e(al_11a7c870[0]),
    .f(al_11a7c870[1]),
    .o(al_3e345b21[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_79894a85 (
    .a(al_ac18355b[4]),
    .b(al_d0a384c4[4]),
    .c(al_1e043bfe[4]),
    .d(al_b0a8403e[4]),
    .e(al_11a7c870[0]),
    .f(al_11a7c870[1]),
    .o(al_3e345b21[4]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    al_7581c23d (
    .a(al_ef78cbcb),
    .b(al_1f97cafb[0]),
    .c(al_1f97cafb[1]),
    .o(al_ba1a11d0));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_2be263e9 (
    .a(al_ba1a11d0),
    .b(al_11a7c870[0]),
    .o(al_1f1dc264[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*~A))"),
    .INIT(8'hb4))
    al_c709433b (
    .a(al_ba1a11d0),
    .b(al_11a7c870[0]),
    .c(al_11a7c870[1]),
    .o(al_1f1dc264[1]));
  AL_MAP_LUT4 #(
    .EQN("(D@(~C*~(B*~A)))"),
    .INIT(16'hf40b))
    al_9c9984e0 (
    .a(al_cefb896),
    .b(al_485702b6),
    .c(al_13f9c71c),
    .d(al_864a13d9[0]),
    .o(al_b528368c[0]));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~C*~(B*~A)))"),
    .INIT(32'hf4ff0b00))
    al_ddc73220 (
    .a(al_cefb896),
    .b(al_485702b6),
    .c(al_13f9c71c),
    .d(al_864a13d9[0]),
    .e(al_864a13d9[1]),
    .o(al_b528368c[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_e1efde68 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_1f1dc264[0]),
    .d(al_1f1dc264[1]),
    .o(al_21302b8a));
  AL_DFF_0 al_a36fbed5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21302b8a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e2903f5));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(C*~A))"),
    .INIT(16'h639c))
    al_8f7e4a98 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_1f1dc264[0]),
    .d(al_1f1dc264[1]),
    .o(al_e1208a36[1]));
  AL_DFF_0 al_f2d0fd5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1208a36[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_79dddfae));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_47fab679 (
    .a(al_864a13d9[0]),
    .b(al_864a13d9[1]),
    .o(al_a83e1130[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(~E*~D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffffffcca0a0a080))
    al_414be30e (
    .a(al_ebb9528c),
    .b(al_ba1a11d0),
    .c(al_a83e1130[0]),
    .d(al_11a7c870[0]),
    .e(al_11a7c870[1]),
    .f(al_413c0926[0]),
    .o(al_6779071c[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_e29bfd1 (
    .a(al_864a13d9[0]),
    .b(al_864a13d9[1]),
    .o(al_a83e1130[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(~E*D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffffccffa0a080a0))
    al_f322d7b2 (
    .a(al_ebb9528c),
    .b(al_ba1a11d0),
    .c(al_a83e1130[1]),
    .d(al_11a7c870[0]),
    .e(al_11a7c870[1]),
    .f(al_413c0926[1]),
    .o(al_6779071c[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d272047f (
    .a(al_864a13d9[0]),
    .b(al_864a13d9[1]),
    .o(al_a83e1130[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(E*~D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffccffffa080a0a0))
    al_62d8706c (
    .a(al_ebb9528c),
    .b(al_ba1a11d0),
    .c(al_a83e1130[2]),
    .d(al_11a7c870[0]),
    .e(al_11a7c870[1]),
    .f(al_413c0926[2]),
    .o(al_6779071c[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_b46faa2b (
    .a(al_864a13d9[0]),
    .b(al_864a13d9[1]),
    .o(al_a83e1130[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    al_26aab38d (
    .a(al_cefb896),
    .b(al_485702b6),
    .c(al_13f9c71c),
    .o(al_ebb9528c));
  AL_MAP_LUT6 #(
    .EQN("(~(E*D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hccffffff80a0a0a0))
    al_102306d (
    .a(al_ebb9528c),
    .b(al_ba1a11d0),
    .c(al_a83e1130[3]),
    .d(al_11a7c870[0]),
    .e(al_11a7c870[1]),
    .f(al_413c0926[3]),
    .o(al_6779071c[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_4b2167ac (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[11]),
    .d(al_e9ebbe15[11]),
    .e(al_c5c971b[11]),
    .f(al_51cc7f19[11]),
    .o(al_55edb257));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_cb49694e (
    .a(al_55edb257),
    .b(al_9e2903f5),
    .c(al_8941a5fb[11]),
    .o(al_e6e3a9da[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_2f6034f7 (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[12]),
    .d(al_e9ebbe15[12]),
    .e(al_c5c971b[12]),
    .f(al_51cc7f19[12]),
    .o(al_7f538ee3));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_d3d65a08 (
    .a(al_7f538ee3),
    .b(al_9e2903f5),
    .c(al_8941a5fb[12]),
    .o(al_e6e3a9da[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_2c7fc870 (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[13]),
    .d(al_e9ebbe15[13]),
    .e(al_c5c971b[13]),
    .f(al_51cc7f19[13]),
    .o(al_c678831f));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_a17d1107 (
    .a(al_c678831f),
    .b(al_9e2903f5),
    .c(al_8941a5fb[13]),
    .o(al_e6e3a9da[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_94835225 (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[14]),
    .d(al_e9ebbe15[14]),
    .e(al_c5c971b[14]),
    .f(al_51cc7f19[14]),
    .o(al_f53b3776));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_7e5255b4 (
    .a(al_f53b3776),
    .b(al_9e2903f5),
    .c(al_8941a5fb[14]),
    .o(al_e6e3a9da[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_3945b9b (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[15]),
    .d(al_e9ebbe15[15]),
    .e(al_c5c971b[15]),
    .f(al_51cc7f19[15]),
    .o(al_1d2d788b));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_8c62db (
    .a(al_1d2d788b),
    .b(al_9e2903f5),
    .c(al_8941a5fb[15]),
    .o(al_e6e3a9da[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_9b15434 (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[16]),
    .d(al_e9ebbe15[16]),
    .e(al_c5c971b[16]),
    .f(al_51cc7f19[16]),
    .o(al_a2fce1));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_cd4f4fdb (
    .a(al_a2fce1),
    .b(al_9e2903f5),
    .c(al_8941a5fb[16]),
    .o(al_e6e3a9da[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_443c4a0e (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[17]),
    .d(al_e9ebbe15[17]),
    .e(al_c5c971b[17]),
    .f(al_51cc7f19[17]),
    .o(al_eb7b08f0));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_29f0e886 (
    .a(al_eb7b08f0),
    .b(al_9e2903f5),
    .c(al_8941a5fb[17]),
    .o(al_e6e3a9da[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_c0c382fe (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[2]),
    .d(al_e9ebbe15[2]),
    .e(al_c5c971b[2]),
    .f(al_51cc7f19[2]),
    .o(al_e355d8ea));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_bcf6c6e5 (
    .a(al_e355d8ea),
    .b(al_9e2903f5),
    .c(al_8941a5fb[2]),
    .o(al_e6e3a9da[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_139350d5 (
    .a(al_c0079c57[0]),
    .b(al_e2c05b54[0]),
    .c(al_a2f64ded[0]),
    .d(al_b1db173b[0]),
    .e(al_f2dedfad[0]),
    .f(al_f2dedfad[1]),
    .o(al_516990df));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_efb4808c (
    .a(al_516990df),
    .b(al_9860067e),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[0]),
    .f(al_75c0d27f[0]),
    .o(al_fcd9679a[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_5ccf9a4f (
    .a(al_fcd9679a[0]),
    .b(al_e2c05b54[0]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_7a57f678[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_b3adeec3 (
    .a(al_fcd9679a[0]),
    .b(al_b1db173b[0]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_73725553[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_f5b0ad2 (
    .a(al_fcd9679a[0]),
    .b(al_a2f64ded[0]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_402dba27[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_5bec6454 (
    .a(al_fcd9679a[0]),
    .b(al_c0079c57[0]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_ff390a8f[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_d983dc9 (
    .a(al_7a57f678[0]),
    .b(al_73725553[0]),
    .c(al_402dba27[0]),
    .d(al_ff390a8f[0]),
    .e(al_864a13d9[0]),
    .f(al_864a13d9[1]),
    .o(al_46448d9c[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_9e158cd5 (
    .a(al_c0079c57[1]),
    .b(al_e2c05b54[1]),
    .c(al_a2f64ded[1]),
    .d(al_b1db173b[1]),
    .e(al_f2dedfad[0]),
    .f(al_f2dedfad[1]),
    .o(al_d87d83a));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'h22222ee2e22eeeee))
    al_b3aadb4e (
    .a(al_d87d83a),
    .b(al_9860067e),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[1]),
    .f(al_75c0d27f[1]),
    .o(al_f16dd8ea));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((~D*C))+~B*A*~((~D*C))+~(~B)*A*(~D*C)+~B*A*(~D*C))"),
    .INIT(16'hcc5c))
    al_2fe8ed0 (
    .a(al_f16dd8ea),
    .b(al_e2c05b54[1]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_7a57f678[1]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((D*C))+~B*A*~((D*C))+~(~B)*A*(D*C)+~B*A*(D*C))"),
    .INIT(16'h5ccc))
    al_6831172c (
    .a(al_f16dd8ea),
    .b(al_b1db173b[1]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_73725553[1]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((D*~C))+~B*A*~((D*~C))+~(~B)*A*(D*~C)+~B*A*(D*~C))"),
    .INIT(16'hc5cc))
    al_624e8802 (
    .a(al_f16dd8ea),
    .b(al_a2f64ded[1]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_402dba27[1]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((~D*~C))+~B*A*~((~D*~C))+~(~B)*A*(~D*~C)+~B*A*(~D*~C))"),
    .INIT(16'hccc5))
    al_b115619b (
    .a(al_f16dd8ea),
    .b(al_c0079c57[1]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_ff390a8f[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_4271df50 (
    .a(al_7a57f678[1]),
    .b(al_73725553[1]),
    .c(al_402dba27[1]),
    .d(al_ff390a8f[1]),
    .e(al_864a13d9[0]),
    .f(al_864a13d9[1]),
    .o(al_46448d9c[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_63e3c27f (
    .a(al_c0079c57[2]),
    .b(al_e2c05b54[2]),
    .c(al_a2f64ded[2]),
    .d(al_b1db173b[2]),
    .e(al_f2dedfad[0]),
    .f(al_f2dedfad[1]),
    .o(al_cb650584));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_34c59877 (
    .a(al_cb650584),
    .b(al_9860067e),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[2]),
    .f(al_75c0d27f[2]),
    .o(al_fcd9679a[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_54731ede (
    .a(al_fcd9679a[2]),
    .b(al_e2c05b54[2]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_7a57f678[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_ae12dc1f (
    .a(al_fcd9679a[2]),
    .b(al_b1db173b[2]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_73725553[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_721ef8db (
    .a(al_fcd9679a[2]),
    .b(al_a2f64ded[2]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_402dba27[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_a8adfcf2 (
    .a(al_fcd9679a[2]),
    .b(al_c0079c57[2]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_ff390a8f[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_455d67aa (
    .a(al_7a57f678[2]),
    .b(al_73725553[2]),
    .c(al_402dba27[2]),
    .d(al_ff390a8f[2]),
    .e(al_864a13d9[0]),
    .f(al_864a13d9[1]),
    .o(al_46448d9c[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_6913513e (
    .a(al_c0079c57[3]),
    .b(al_e2c05b54[3]),
    .c(al_a2f64ded[3]),
    .d(al_b1db173b[3]),
    .e(al_f2dedfad[0]),
    .f(al_f2dedfad[1]),
    .o(al_254e8e6));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_e32ca926 (
    .a(al_254e8e6),
    .b(al_9860067e),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[3]),
    .f(al_75c0d27f[3]),
    .o(al_fcd9679a[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_29eed166 (
    .a(al_fcd9679a[3]),
    .b(al_e2c05b54[3]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_7a57f678[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_768cf200 (
    .a(al_fcd9679a[3]),
    .b(al_b1db173b[3]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_73725553[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_5895f0b4 (
    .a(al_fcd9679a[3]),
    .b(al_a2f64ded[3]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_402dba27[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_daf6b121 (
    .a(al_fcd9679a[3]),
    .b(al_c0079c57[3]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_ff390a8f[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_6f4b54a4 (
    .a(al_7a57f678[3]),
    .b(al_73725553[3]),
    .c(al_402dba27[3]),
    .d(al_ff390a8f[3]),
    .e(al_864a13d9[0]),
    .f(al_864a13d9[1]),
    .o(al_46448d9c[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_1ae7908b (
    .a(al_c0079c57[4]),
    .b(al_e2c05b54[4]),
    .c(al_a2f64ded[4]),
    .d(al_b1db173b[4]),
    .e(al_f2dedfad[0]),
    .f(al_f2dedfad[1]),
    .o(al_1dde650a));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*(D@C)))*~(B)+~A*(E*(D@C))*~(B)+~(~A)*(E*(D@C))*B+~A*(E*(D@C))*B)"),
    .INIT(32'h1dd11111))
    al_798d54e9 (
    .a(al_1dde650a),
    .b(al_9860067e),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[4]),
    .o(al_fcd9679a[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_352be493 (
    .a(al_fcd9679a[4]),
    .b(al_e2c05b54[4]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_7a57f678[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_e6852db6 (
    .a(al_fcd9679a[4]),
    .b(al_b1db173b[4]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_73725553[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_6185bb3b (
    .a(al_fcd9679a[4]),
    .b(al_a2f64ded[4]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_402dba27[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_fabb67ad (
    .a(al_fcd9679a[4]),
    .b(al_c0079c57[4]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_ff390a8f[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_4940f80c (
    .a(al_7a57f678[4]),
    .b(al_73725553[4]),
    .c(al_402dba27[4]),
    .d(al_ff390a8f[4]),
    .e(al_864a13d9[0]),
    .f(al_864a13d9[1]),
    .o(al_46448d9c[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_4739feb7 (
    .a(al_6860fc86),
    .b(al_74055ffa),
    .c(al_7b43c1e),
    .d(al_8cddf958),
    .o(al_221aa358));
  AL_MAP_LUT6 #(
    .EQN("(F*~(~E*~D*C*~B*A))"),
    .INIT(64'hffffffdf00000000))
    al_fbf79e64 (
    .a(al_94f083a0),
    .b(al_a0789cd8),
    .c(al_c711503f),
    .d(al_cfa51fb3[0]),
    .e(al_cfa51fb3[1]),
    .f(al_6dee9bef),
    .o(al_50105215));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    al_22504ba4 (
    .a(al_221aa358),
    .b(al_2dc3e45),
    .c(al_50105215),
    .o(al_16929b7c[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    al_56eca0d8 (
    .a(al_221aa358),
    .b(al_f027c275),
    .c(al_369e229d[0]),
    .o(al_63714fc7));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*B*~(E*A)))"),
    .INIT(32'h00bf003f))
    al_aa246cc3 (
    .a(al_79dddfae),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_369e229d[2]),
    .e(al_c360bf4c[2]),
    .o(al_6d69b644));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E*~(~D*~(B*~A))))"),
    .INIT(32'h000b0f0f))
    al_5ac51d26 (
    .a(al_16929b7c[0]),
    .b(al_63714fc7),
    .c(al_86941e27),
    .d(al_4eef0b42),
    .e(al_6d69b644),
    .o(al_edda145c[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_d4f8d4a7 (
    .a(al_ca418906),
    .b(al_a0789cd8),
    .c(al_c711503f),
    .o(al_2dc3e45));
  AL_MAP_LUT4 #(
    .EQN("(A*(~(B)*~(C)*~(D)+B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D+~(B)*C*D))"),
    .INIT(16'h282a))
    al_41aa7f30 (
    .a(al_13f9c71c),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_f7e9a10b),
    .o(al_86941e27));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~(~D*~(C*~(F*~(B*~A)))))"),
    .INIT(64'hffff00bfffff000f))
    al_a8eb22a1 (
    .a(al_58fb4752[3]),
    .b(al_58fb4752[4]),
    .c(al_f7a41bbb),
    .d(al_369e229d[0]),
    .e(al_369e229d[1]),
    .f(al_ad9637b9),
    .o(al_4eef0b42));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_caf162e4 (
    .a(al_6896ad14),
    .b(al_ad9637b9),
    .o(al_6dee9bef));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d36fe55e (
    .a(al_221aa358),
    .b(al_2dc3e45),
    .o(al_9d2235cc));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(E*~((D*~A))*~(B)+E*(D*~A)*~(B)+~(E)*(D*~A)*B+E*(D*~A)*B))"),
    .INIT(32'h7f3f4f0f))
    al_3ea12990 (
    .a(al_79dddfae),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_c360bf4c[2]),
    .e(al_165f2734),
    .o(al_81850512));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1c1f))
    al_5e320807 (
    .a(al_79dddfae),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_f7e9a10b),
    .o(al_1d4e62f6));
  AL_MAP_LUT6 #(
    .EQN("~((C*~(E*~(~B*~A)))*~(D)*~(F)+(C*~(E*~(~B*~A)))*D*~(F)+~((C*~(E*~(~B*~A))))*D*F+(C*~(E*~(~B*~A)))*D*F)"),
    .INIT(64'h00ff00ffefef0f0f))
    al_5cfd5fc9 (
    .a(al_9d2235cc),
    .b(al_114b0fe8),
    .c(al_81850512),
    .d(al_1d4e62f6),
    .e(al_6ad3f77e),
    .f(al_369e229d[2]),
    .o(al_edda145c[1]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    al_edd1c7a1 (
    .a(al_79dddfae),
    .b(al_369e229d[0]),
    .c(al_c360bf4c[2]),
    .d(al_165f2734),
    .o(al_1af39dee));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfcf05500fcff5500))
    al_70fe5a6c (
    .a(al_1af39dee),
    .b(al_79dddfae),
    .c(al_369e229d[0]),
    .d(al_369e229d[1]),
    .e(al_369e229d[2]),
    .f(al_f7e9a10b),
    .o(al_edda145c[2]));
  AL_MAP_LUT5 #(
    .EQN("((~B*A)*~(C)*~(D)*~(E)+(~B*A)*C*~(D)*~(E)+~((~B*A))*~(C)*D*~(E)+(~B*A)*~(C)*D*~(E)+~((~B*A))*C*~(D)*E+(~B*A)*C*~(D)*E+~((~B*A))*~(C)*D*E+(~B*A)*~(C)*D*E+~((~B*A))*C*D*E+(~B*A)*C*D*E)"),
    .INIT(32'hfff00f22))
    al_5bf0d77 (
    .a(al_85567015),
    .b(al_b3701730),
    .c(al_ef78cbcb),
    .d(al_1f97cafb[0]),
    .e(al_1f97cafb[1]),
    .o(al_9adc03c8[0]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(~C*B*A))"),
    .INIT(16'hff08))
    al_15956b40 (
    .a(al_85567015),
    .b(al_b3701730),
    .c(al_1f97cafb[0]),
    .d(al_1f97cafb[1]),
    .o(al_9adc03c8[1]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_e3337a5d (
    .a(al_1c962936),
    .b(al_77041990),
    .c(al_31da793),
    .o(al_3a754a7b));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_20ace8ce (
    .a(al_c72051a5),
    .b(al_77041990),
    .c(al_31da793),
    .o(al_2e8f51d8));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_412875c7 (
    .a(al_1316088),
    .b(al_77041990),
    .c(al_31da793),
    .o(al_e82b7392));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_56cdacf (
    .a(al_cf11b78b[2]),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_369e229d[2]),
    .e(al_898823b1),
    .o(al_77041990));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_56f8a75 (
    .a(al_d8e50712),
    .b(al_77041990),
    .c(al_31da793),
    .o(al_7326000a));
  AL_DFF_0 al_a2f96b64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ddeaf309),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_4135f4fc));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    al_e740e7a1 (
    .a(al_7c6fd728),
    .b(al_4135f4fc),
    .c(al_165f2734),
    .o(al_ddeaf309));
  AL_DFF_0 al_e72a4c1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21bd4e5d[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_1d36bc6d));
  AL_DFF_0 al_17964f7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21bd4e5d[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_b0fb8887));
  AL_DFF_0 al_ff7298e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21bd4e5d[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_a9552c76));
  AL_DFF_0 al_6ef6f503 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21bd4e5d[3]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_4331638));
  AL_DFF_0 al_d349a677 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21bd4e5d[4]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2a6634d6));
  AL_DFF_0 al_de6092fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6824a1b1[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_c54166ab));
  AL_DFF_0 al_396fada (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6824a1b1[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_41e1e6ea));
  AL_DFF_0 al_1f0306f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6824a1b1[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_a01620de));
  AL_DFF_0 al_e9b4eddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6824a1b1[3]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_27a9ba79));
  AL_DFF_0 al_8bf78f82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6d285e98[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e59c045a));
  AL_DFF_0 al_a93c35dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6d285e98[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_41fff7fc));
  AL_DFF_0 al_4145b995 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6d285e98[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2acc39d8));
  AL_DFF_0 al_6a0840c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6d285e98[3]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_27a5f0e3));
  AL_DFF_0 al_8c5008ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_579d2a90[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_dc7ca9c3));
  AL_DFF_0 al_f854996d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_579d2a90[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_3b67e711));
  AL_DFF_0 al_f4f65b50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_579d2a90[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_764705a7));
  AL_DFF_0 al_97382205 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_579d2a90[3]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e9b4dc12));
  AL_DFF_0 al_3b17dd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2f1f444b[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_fa80f9c4));
  AL_DFF_0 al_da5b78c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2f1f444b[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_65940b21));
  AL_DFF_0 al_94ea8dfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2f1f444b[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e5dd3f8d));
  AL_DFF_0 al_bfc22ae5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2f1f444b[3]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_749a40e9));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_e156b03f (
    .a(al_369e229d[0]),
    .b(al_369e229d[1]),
    .c(al_369e229d[2]),
    .o(al_19014a7b));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_c8c492a5 (
    .a(al_19014a7b),
    .b(al_8941a5fb[0]),
    .c(al_8941a5fb[1]),
    .o(al_c72051a5));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_160f6acd (
    .a(al_c72051a5),
    .b(al_c360bf4c[2]),
    .o(al_32770943));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_2ff73ade (
    .a(al_32770943),
    .b(al_e59c045a),
    .c(al_41fff7fc),
    .d(al_2acc39d8),
    .e(al_27a5f0e3),
    .f(al_c74d7793),
    .o(al_6d285e98[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_10ece330 (
    .a(al_32770943),
    .b(al_e59c045a),
    .c(al_c74d7793),
    .o(al_6d285e98[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_517d67b7 (
    .a(al_32770943),
    .b(al_e59c045a),
    .c(al_41fff7fc),
    .d(al_c74d7793),
    .o(al_6d285e98[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_36ad524f (
    .a(al_32770943),
    .b(al_e59c045a),
    .c(al_41fff7fc),
    .d(al_2acc39d8),
    .e(al_c74d7793),
    .o(al_6d285e98[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_83503389 (
    .a(al_19014a7b),
    .b(al_8941a5fb[0]),
    .c(al_8941a5fb[1]),
    .o(al_1316088));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_e639f921 (
    .a(al_1316088),
    .b(al_c360bf4c[2]),
    .o(al_f01cf98));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_a710c197 (
    .a(al_f01cf98),
    .b(al_dc7ca9c3),
    .c(al_3b67e711),
    .d(al_764705a7),
    .e(al_e9b4dc12),
    .f(al_82bb1e86),
    .o(al_579d2a90[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_8a0e0863 (
    .a(al_f01cf98),
    .b(al_dc7ca9c3),
    .c(al_82bb1e86),
    .o(al_579d2a90[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_7a5c42ca (
    .a(al_f01cf98),
    .b(al_dc7ca9c3),
    .c(al_3b67e711),
    .d(al_82bb1e86),
    .o(al_579d2a90[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_1c0a6c46 (
    .a(al_f01cf98),
    .b(al_dc7ca9c3),
    .c(al_3b67e711),
    .d(al_764705a7),
    .e(al_82bb1e86),
    .o(al_579d2a90[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_897a5815 (
    .a(al_19014a7b),
    .b(al_8941a5fb[0]),
    .c(al_8941a5fb[1]),
    .o(al_d8e50712));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9da2f175 (
    .a(al_d8e50712),
    .b(al_c360bf4c[2]),
    .o(al_22cea9d));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_442f0d33 (
    .a(al_22cea9d),
    .b(al_fa80f9c4),
    .c(al_65940b21),
    .d(al_e5dd3f8d),
    .e(al_749a40e9),
    .f(al_3b347f86),
    .o(al_2f1f444b[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_24afdc66 (
    .a(al_22cea9d),
    .b(al_fa80f9c4),
    .c(al_3b347f86),
    .o(al_2f1f444b[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_50cc8729 (
    .a(al_22cea9d),
    .b(al_fa80f9c4),
    .c(al_65940b21),
    .d(al_3b347f86),
    .o(al_2f1f444b[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_a06d36c5 (
    .a(al_22cea9d),
    .b(al_fa80f9c4),
    .c(al_65940b21),
    .d(al_e5dd3f8d),
    .e(al_3b347f86),
    .o(al_2f1f444b[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_83b6ca34 (
    .a(al_19014a7b),
    .b(al_8941a5fb[0]),
    .c(al_8941a5fb[1]),
    .o(al_1c962936));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_121da31c (
    .a(al_1c962936),
    .b(al_c360bf4c[2]),
    .o(al_f7f8cb1));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_dcca4fc (
    .a(al_f7f8cb1),
    .b(al_c54166ab),
    .c(al_41e1e6ea),
    .d(al_a01620de),
    .e(al_27a9ba79),
    .f(al_1cf815c1),
    .o(al_6824a1b1[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_c9204305 (
    .a(al_f7f8cb1),
    .b(al_c54166ab),
    .c(al_1cf815c1),
    .o(al_6824a1b1[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_721f6127 (
    .a(al_f7f8cb1),
    .b(al_c54166ab),
    .c(al_41e1e6ea),
    .d(al_1cf815c1),
    .o(al_6824a1b1[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_63012592 (
    .a(al_f7f8cb1),
    .b(al_c54166ab),
    .c(al_41e1e6ea),
    .d(al_a01620de),
    .e(al_1cf815c1),
    .o(al_6824a1b1[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_880e1570 (
    .a(al_6d285e98[3]),
    .b(al_6d285e98[0]),
    .c(al_6d285e98[1]),
    .d(al_6d285e98[2]),
    .o(al_86261d41[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_9bec58a7 (
    .a(al_579d2a90[3]),
    .b(al_579d2a90[0]),
    .c(al_579d2a90[1]),
    .d(al_579d2a90[2]),
    .o(al_86261d41[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_b548977 (
    .a(al_2f1f444b[3]),
    .b(al_2f1f444b[0]),
    .c(al_2f1f444b[1]),
    .d(al_2f1f444b[2]),
    .o(al_86261d41[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_eb8c44ab (
    .a(al_6824a1b1[3]),
    .b(al_6824a1b1[0]),
    .c(al_6824a1b1[1]),
    .d(al_6824a1b1[2]),
    .o(al_86261d41[0]));
  AL_DFF_0 al_af83d51b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_86261d41[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cf815c1));
  AL_DFF_0 al_5b04d785 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_86261d41[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c74d7793));
  AL_DFF_0 al_5bc607d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_86261d41[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82bb1e86));
  AL_DFF_0 al_7d427b78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_86261d41[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b347f86));
  AL_DFF_0 al_162ed9d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7ab735a9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_833f5c05));
  AL_DFF_0 al_77a1dcc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[24]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e707cc02));
  AL_DFF_0 al_1a78b677 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[25]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_464fb058));
  AL_DFF_0 al_d4e3f545 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[26]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_9d701591));
  AL_DFF_0 al_1dbdd7a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[27]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_b1edca88));
  AL_DFF_0 al_11daf923 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[28]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_48aee091));
  AL_DFF_0 al_a12f7e4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[29]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_3185ed47));
  AL_DFF_0 al_ea6bea1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[30]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2e96480));
  AL_DFF_0 al_ae914b7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[31]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_9264d6ce));
  AL_DFF_0 al_d1cfa2ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[32]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e2bcb10));
  AL_DFF_0 al_83e3b56c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[33]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_1b6a0af9));
  AL_DFF_0 al_472e0c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[34]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_5d3dfa86));
  AL_DFF_0 al_3f627349 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[35]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_403fbf52));
  AL_DFF_0 al_eb2fb067 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[36]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_8287cea7));
  AL_DFF_0 al_ec4c5bfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[37]),
    .en(al_3a754a7b),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_a4914504));
  AL_DFF_0 al_b7ceb988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_37a27dff),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3df83ccd));
  AL_DFF_0 al_d4c824f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[24]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e2740cd5));
  AL_DFF_0 al_83f5c8fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[25]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_fd5ac0c0));
  AL_DFF_0 al_3185a856 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[26]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_bd5f3c97));
  AL_DFF_0 al_5fe65d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[27]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_364b2d93));
  AL_DFF_0 al_13bdc847 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[28]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_10d1f7da));
  AL_DFF_0 al_cdc30aff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[29]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_bfe0071c));
  AL_DFF_0 al_66821e2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[30]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_22a3e261));
  AL_DFF_0 al_314169ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[31]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_9dee74a8));
  AL_DFF_0 al_47c9e798 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[32]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_25de7719));
  AL_DFF_0 al_6bf8e393 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[33]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_6a2ba50d));
  AL_DFF_0 al_f66cbd8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[34]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_55c1f3f8));
  AL_DFF_0 al_333fd08c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[35]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_53439d34));
  AL_DFF_0 al_31e1c929 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[36]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_dedd5989));
  AL_DFF_0 al_6fbdb1d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[37]),
    .en(al_2e8f51d8),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_a1d2ac98));
  AL_DFF_0 al_8b7f22d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d1dcebd4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_61792012));
  AL_DFF_0 al_8a418ffc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[24]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_4743871));
  AL_DFF_0 al_fd05b2ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[25]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_6bbd7053));
  AL_DFF_0 al_2eaf3d47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[26]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e4c2295a));
  AL_DFF_0 al_366b2b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[27]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_28da8a0d));
  AL_DFF_0 al_23dc90c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[28]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_539c7732));
  AL_DFF_0 al_5f3100c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[29]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_6692b66c));
  AL_DFF_0 al_33eb907 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[30]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_3647cd0));
  AL_DFF_0 al_4fd312b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[31]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_b62c6ace));
  AL_DFF_0 al_b3e16e72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[32]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_49d43cfa));
  AL_DFF_0 al_8b03ba95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[33]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_c32d8f29));
  AL_DFF_0 al_b5154dd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[34]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2f5e01b7));
  AL_DFF_0 al_584c3e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[35]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2a5fa8c));
  AL_DFF_0 al_703dd454 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[36]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_b4d9e182));
  AL_DFF_0 al_70e1b2ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[37]),
    .en(al_e82b7392),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_34ff0ff5));
  AL_DFF_0 al_d1acce72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3303cc51),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_286587c2));
  AL_DFF_0 al_75c6b3d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[24]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f498aaed));
  AL_DFF_0 al_fcc36f01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[25]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_dd9df6a3));
  AL_DFF_0 al_d01c1a17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[26]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_26b95353));
  AL_DFF_0 al_661c50f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[27]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e1521e17));
  AL_DFF_0 al_5bc73f38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[28]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_a448873e));
  AL_DFF_0 al_81986860 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[29]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e80539a7));
  AL_DFF_0 al_4b3dd6b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[30]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_9526df3b));
  AL_DFF_0 al_3de56ac7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[31]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_c959a932));
  AL_DFF_0 al_d5e611ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[32]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_fc1936a5));
  AL_DFF_0 al_b22badde (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[33]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_66bed231));
  AL_DFF_0 al_3c848e8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[34]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_a04a63d4));
  AL_DFF_0 al_52bf08b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[35]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_ebe69372));
  AL_DFF_0 al_386aaffe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[36]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_e0a71537));
  AL_DFF_0 al_36fc2de6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[37]),
    .en(al_7326000a),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_18d4d578));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_8911ed6b (
    .a(al_c72051a5),
    .b(al_77041990),
    .c(al_3df83ccd),
    .d(al_31da793),
    .e(al_cbaa3056),
    .o(al_37a27dff));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_dd1adb06 (
    .a(al_1c962936),
    .b(al_77041990),
    .c(al_833f5c05),
    .d(al_31da793),
    .e(al_cbaa3056),
    .o(al_7ab735a9));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_a265ca7b (
    .a(al_d8e50712),
    .b(al_77041990),
    .c(al_286587c2),
    .d(al_31da793),
    .e(al_cbaa3056),
    .o(al_3303cc51));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_100b46fb (
    .a(al_1316088),
    .b(al_77041990),
    .c(al_61792012),
    .d(al_31da793),
    .e(al_cbaa3056),
    .o(al_d1dcebd4));
  AL_DFF_0 al_58df8c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4bc24ece[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_31da793));
  AL_DFF_0 al_f9e101ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_61614b33[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_19e106e3));
  AL_DFF_0 al_bb1b8548 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d6f3e78f),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_a70d3eb4));
  AL_MAP_LUT6 #(
    .EQN("(~C*~(~D*~(~F*~E*B*A)))"),
    .INIT(64'h0f000f000f000f08))
    al_91b6f3c0 (
    .a(al_85567015),
    .b(al_732fadca),
    .c(al_ef78cbcb),
    .d(al_a70d3eb4),
    .e(al_1f97cafb[0]),
    .f(al_1f97cafb[1]),
    .o(al_d6f3e78f));
  AL_DFF_0 al_7ed97c68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a77bd6b4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf11b78b[2]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_3b62477c (
    .a(al_6896ad14),
    .b(al_9e2903f5),
    .c(al_369e229d[0]),
    .d(al_369e229d[1]),
    .e(al_369e229d[2]),
    .o(al_a77bd6b4));
  AL_DFF_0 al_8d8364d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eae09b27),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbeafa67[4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    al_cac4ae0b (
    .a(al_7c6fd728),
    .b(al_cbeafa67[4]),
    .c(al_8941a5fb[2]),
    .d(al_cbaa3056),
    .o(al_eae09b27));
  AL_DFF_0 al_8656e7ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_aaf3456[0]));
  AL_DFF_0 al_54cc5d0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_aaf3456[1]));
  AL_DFF_0 al_19a8a26c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_d76fa964[4]));
  AL_DFF_0 al_ecd27a70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_edda145c[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_369e229d[0]));
  AL_DFF_0 al_4fa1cac9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_edda145c[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_369e229d[1]));
  AL_DFF_0 al_f83c3214 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_edda145c[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_369e229d[2]));
  AL_DFF_0 al_14761d07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9adc03c8[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_1f97cafb[0]));
  AL_DFF_0 al_38665934 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9adc03c8[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_1f97cafb[1]));
  AL_DFF_0 al_c985b016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff390a8f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0079c57[0]));
  AL_DFF_0 al_5acc339e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff390a8f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0079c57[1]));
  AL_DFF_0 al_32bafbce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff390a8f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0079c57[2]));
  AL_DFF_0 al_76f2fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff390a8f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0079c57[3]));
  AL_DFF_0 al_afd950e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff390a8f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0079c57[4]));
  AL_DFF_0 al_349e0416 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7a57f678[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e2c05b54[0]));
  AL_DFF_0 al_1eee66f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7a57f678[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e2c05b54[1]));
  AL_DFF_0 al_cbc71ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7a57f678[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e2c05b54[2]));
  AL_DFF_0 al_9e2c88ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7a57f678[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e2c05b54[3]));
  AL_DFF_0 al_43701ca2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7a57f678[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e2c05b54[4]));
  AL_DFF_0 al_4981eda (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_402dba27[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a2f64ded[0]));
  AL_DFF_0 al_74c16ea8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_402dba27[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a2f64ded[1]));
  AL_DFF_0 al_17ed7ae0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_402dba27[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a2f64ded[2]));
  AL_DFF_0 al_e454f1c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_402dba27[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a2f64ded[3]));
  AL_DFF_0 al_ef9a182a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_402dba27[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a2f64ded[4]));
  AL_DFF_0 al_91af0c6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_73725553[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1db173b[0]));
  AL_DFF_0 al_91c6fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_73725553[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1db173b[1]));
  AL_DFF_0 al_fd7d698c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_73725553[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1db173b[2]));
  AL_DFF_0 al_50f58047 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_73725553[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1db173b[3]));
  AL_DFF_0 al_6bb197db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_73725553[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b1db173b[4]));
  AL_DFF_0 al_701ab94d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e048ecc8[3]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_7fb24d41[3]));
  AL_DFF_0 al_35ff1573 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e048ecc8[4]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_7fb24d41[4]));
  AL_DFF_0 al_af7bd144 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e048ecc8[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_7fb24d41[0]));
  AL_DFF_0 al_a584dcbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e048ecc8[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_7fb24d41[1]));
  AL_DFF_0 al_a0c1c5ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e048ecc8[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_7fb24d41[2]));
  AL_DFF_0 al_8f1730a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[0]));
  AL_DFF_0 al_fc93d5ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[1]));
  AL_DFF_0 al_f9c3a10b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[2]));
  AL_DFF_0 al_4ed1241d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[11]));
  AL_DFF_0 al_a11740f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[12]));
  AL_DFF_0 al_26a4a6d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[13]));
  AL_DFF_0 al_60e9f05e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[14]));
  AL_DFF_0 al_bcbc5f4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[15]));
  AL_DFF_0 al_88322277 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[16]));
  AL_DFF_0 al_e5147979 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[17]));
  AL_DFF_0 al_96214e2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[24]));
  AL_DFF_0 al_ce38f96d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[25]));
  AL_DFF_0 al_d4b0057f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[26]));
  AL_DFF_0 al_1c5fb187 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[27]));
  AL_DFF_0 al_ecb49683 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[28]));
  AL_DFF_0 al_9c7e8211 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[29]));
  AL_DFF_0 al_551cc832 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[30]));
  AL_DFF_0 al_552a9334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[31]));
  AL_DFF_0 al_4170ee51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[32]));
  AL_DFF_0 al_640cd898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[33]));
  AL_DFF_0 al_7b633708 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[34]));
  AL_DFF_0 al_c2d3d617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[35]));
  AL_DFF_0 al_76911a91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[36]));
  AL_DFF_0 al_d42bb655 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[37]));
  AL_DFF_0 al_975c4e2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[44]));
  AL_DFF_0 al_ffad98bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[45]));
  AL_DFF_0 al_909ef30c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc0d6480[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8941a5fb[46]));
  AL_DFF_0 al_ce9a70f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[0]));
  AL_DFF_0 al_5b5d990 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[1]));
  AL_DFF_0 al_d5ab9e59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[2]));
  AL_DFF_0 al_ff9f8409 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[11]));
  AL_DFF_0 al_4ac4bcf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[12]));
  AL_DFF_0 al_924292e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[13]));
  AL_DFF_0 al_4303376a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[14]));
  AL_DFF_0 al_7f9d262e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[15]));
  AL_DFF_0 al_43a1d69f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[16]));
  AL_DFF_0 al_e933e0a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[17]));
  AL_DFF_0 al_efd8d0ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[24]));
  AL_DFF_0 al_934a73e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[25]));
  AL_DFF_0 al_89d1d290 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[26]));
  AL_DFF_0 al_78ec85c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[27]));
  AL_DFF_0 al_590cf679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[28]));
  AL_DFF_0 al_b6802f8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[29]));
  AL_DFF_0 al_2730f170 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[30]));
  AL_DFF_0 al_8fcb6e6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[31]));
  AL_DFF_0 al_b425ca88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[32]));
  AL_DFF_0 al_924db4f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[33]));
  AL_DFF_0 al_846805a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[34]));
  AL_DFF_0 al_be0dac40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[35]));
  AL_DFF_0 al_6fef683f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[36]));
  AL_DFF_0 al_4db4bd40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[37]));
  AL_DFF_0 al_745417b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[44]));
  AL_DFF_0 al_d5e0641b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[45]));
  AL_DFF_0 al_16dc0478 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_ef92c438[0]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_31adc4ab[46]));
  AL_DFF_0 al_25b2d1ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[0]));
  AL_DFF_0 al_9f08ed63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[1]));
  AL_DFF_0 al_b5777354 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[2]));
  AL_DFF_0 al_755c7499 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[11]));
  AL_DFF_0 al_74764c85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[12]));
  AL_DFF_0 al_8738d5f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[13]));
  AL_DFF_0 al_7801c3c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[14]));
  AL_DFF_0 al_b69094d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[15]));
  AL_DFF_0 al_547dd6c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[16]));
  AL_DFF_0 al_5794984b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[17]));
  AL_DFF_0 al_4cbd9f51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[24]));
  AL_DFF_0 al_d7e20414 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[25]));
  AL_DFF_0 al_2d9effa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[26]));
  AL_DFF_0 al_d0229385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[27]));
  AL_DFF_0 al_e50a281c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[28]));
  AL_DFF_0 al_e8ac347c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[29]));
  AL_DFF_0 al_ccf567e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[30]));
  AL_DFF_0 al_898ae1c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[31]));
  AL_DFF_0 al_2093a758 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[32]));
  AL_DFF_0 al_4c7a7572 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[33]));
  AL_DFF_0 al_60bfa78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[34]));
  AL_DFF_0 al_372372f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[35]));
  AL_DFF_0 al_98fc5f25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[36]));
  AL_DFF_0 al_db797196 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[37]));
  AL_DFF_0 al_281f2471 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[44]));
  AL_DFF_0 al_ed9edf48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[45]));
  AL_DFF_0 al_99c4c715 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_ef92c438[1]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_39d4ac28[46]));
  AL_DFF_0 al_df622221 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[0]));
  AL_DFF_0 al_f425d586 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[1]));
  AL_DFF_0 al_c43edca8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[2]));
  AL_DFF_0 al_724e44e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[11]));
  AL_DFF_0 al_56f5f6ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[12]));
  AL_DFF_0 al_250cac37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[13]));
  AL_DFF_0 al_961c648c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[14]));
  AL_DFF_0 al_ad84d3d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[15]));
  AL_DFF_0 al_f167b47d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[16]));
  AL_DFF_0 al_fa0bc38d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[17]));
  AL_DFF_0 al_8871f500 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[24]));
  AL_DFF_0 al_858e2717 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[25]));
  AL_DFF_0 al_e5e3c355 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[26]));
  AL_DFF_0 al_4831791a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[27]));
  AL_DFF_0 al_c357a2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[28]));
  AL_DFF_0 al_a6e19028 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[29]));
  AL_DFF_0 al_ffa9b04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[30]));
  AL_DFF_0 al_9f215b99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[31]));
  AL_DFF_0 al_96ca3163 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[32]));
  AL_DFF_0 al_866ecfe2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[33]));
  AL_DFF_0 al_97a3f560 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[34]));
  AL_DFF_0 al_588995ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[35]));
  AL_DFF_0 al_c192c7f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[36]));
  AL_DFF_0 al_73557936 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[37]));
  AL_DFF_0 al_21b16be7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[44]));
  AL_DFF_0 al_9a59907c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[45]));
  AL_DFF_0 al_efd47c9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_ef92c438[2]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2697e1b1[46]));
  AL_DFF_0 al_534a69e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[0]));
  AL_DFF_0 al_ef5802f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[1]));
  AL_DFF_0 al_90ac57d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[2]));
  AL_DFF_0 al_80c6bd3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[11]));
  AL_DFF_0 al_e11e78c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[12]));
  AL_DFF_0 al_436afcf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[13]));
  AL_DFF_0 al_bac48767 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[14]));
  AL_DFF_0 al_8eda0f22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[15]));
  AL_DFF_0 al_d878fbae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[16]));
  AL_DFF_0 al_e1fe897a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[17]));
  AL_DFF_0 al_bbd43f66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[24]));
  AL_DFF_0 al_44d61045 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[25]));
  AL_DFF_0 al_528b39c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[26]));
  AL_DFF_0 al_ae0b518c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[27]));
  AL_DFF_0 al_c74525c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[28]));
  AL_DFF_0 al_5d958362 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[29]));
  AL_DFF_0 al_fb32cd56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[30]));
  AL_DFF_0 al_8291b2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[31]));
  AL_DFF_0 al_6fec9678 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[32]));
  AL_DFF_0 al_479db912 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[33]));
  AL_DFF_0 al_287c69e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[34]));
  AL_DFF_0 al_c979fe9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[35]));
  AL_DFF_0 al_e68ea7aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[36]));
  AL_DFF_0 al_9090681e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[37]));
  AL_DFF_0 al_5da1fa86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[44]));
  AL_DFF_0 al_4bc6a900 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[45]));
  AL_DFF_0 al_bd0f675 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_ef92c438[3]),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f0541159[46]));
  AL_DFF_0 al_1fa1c699 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b528368c[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_864a13d9[0]));
  AL_DFF_0 al_2f0ae136 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b528368c[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_864a13d9[1]));
  AL_DFF_0 al_dc30b9ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ca7553ae[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f2dedfad[0]));
  AL_DFF_0 al_c7ea1a27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ca7553ae[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f2dedfad[1]));
  AL_DFF_0 al_9477af65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[0]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac18355b[0]));
  AL_DFF_0 al_9ca2b81e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[1]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac18355b[1]));
  AL_DFF_0 al_c4486081 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[2]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac18355b[2]));
  AL_DFF_0 al_c5d92c81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[3]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac18355b[3]));
  AL_DFF_0 al_ca66c89b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[4]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac18355b[4]));
  AL_DFF_0 al_e484c29e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[0]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d0a384c4[0]));
  AL_DFF_0 al_dad1f45e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[1]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d0a384c4[1]));
  AL_DFF_0 al_d06b63e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[2]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d0a384c4[2]));
  AL_DFF_0 al_4379f093 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[3]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d0a384c4[3]));
  AL_DFF_0 al_36c3a592 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[4]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d0a384c4[4]));
  AL_DFF_0 al_8bb0956e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[0]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e043bfe[0]));
  AL_DFF_0 al_22f4af2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[1]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e043bfe[1]));
  AL_DFF_0 al_aa3a0f6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[2]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e043bfe[2]));
  AL_DFF_0 al_17e4cfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[3]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e043bfe[3]));
  AL_DFF_0 al_fc32056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[4]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e043bfe[4]));
  AL_DFF_0 al_f4b3c48a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[0]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0a8403e[0]));
  AL_DFF_0 al_30a155d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[1]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0a8403e[1]));
  AL_DFF_0 al_815d2973 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[2]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0a8403e[2]));
  AL_DFF_0 al_b60b434e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[3]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0a8403e[3]));
  AL_DFF_0 al_17abffab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46448d9c[4]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0a8403e[4]));
  AL_DFF_0 al_879b0e61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f1dc264[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_11a7c870[0]));
  AL_DFF_0 al_81610d72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f1dc264[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_11a7c870[1]));
  AL_DFF_0 al_647bc239 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6779071c[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_413c0926[0]));
  AL_DFF_0 al_ed8ab0c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6779071c[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_413c0926[1]));
  AL_DFF_0 al_b009af3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6779071c[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_413c0926[2]));
  AL_DFF_0 al_4ca95f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6779071c[3]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_413c0926[3]));
  AL_DFF_0 al_37876f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[0]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[0]));
  AL_DFF_0 al_e74fdad9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[1]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[1]));
  AL_DFF_0 al_c8a46844 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[2]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[2]));
  AL_DFF_0 al_5ca7c390 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[11]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[11]));
  AL_DFF_0 al_ef7ffdd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[12]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[12]));
  AL_DFF_0 al_486e4d96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[13]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[13]));
  AL_DFF_0 al_6d4e7a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[14]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[14]));
  AL_DFF_0 al_b7d3832a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[15]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[15]));
  AL_DFF_0 al_c6cb8ccd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[16]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[16]));
  AL_DFF_0 al_b7ac9166 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[17]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[17]));
  AL_DFF_0 al_2fec3957 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[44]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[44]));
  AL_DFF_0 al_ca2bdb07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[45]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[45]));
  AL_DFF_0 al_b14f044f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[46]),
    .en(al_a83e1130[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59b0cd05[46]));
  AL_DFF_0 al_c38ca2fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[0]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[0]));
  AL_DFF_0 al_7d986244 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[1]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[1]));
  AL_DFF_0 al_9dd2d203 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[2]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[2]));
  AL_DFF_0 al_82a999ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[11]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[11]));
  AL_DFF_0 al_76d612a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[12]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[12]));
  AL_DFF_0 al_98f8090e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[13]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[13]));
  AL_DFF_0 al_fa7b684d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[14]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[14]));
  AL_DFF_0 al_6ed9035 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[15]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[15]));
  AL_DFF_0 al_ee5e0940 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[16]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[16]));
  AL_DFF_0 al_6022daae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[17]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[17]));
  AL_DFF_0 al_447bf146 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[44]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[44]));
  AL_DFF_0 al_5095f3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[45]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[45]));
  AL_DFF_0 al_391473ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[46]),
    .en(al_a83e1130[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9ebbe15[46]));
  AL_DFF_0 al_cb8a8e77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[0]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[0]));
  AL_DFF_0 al_a3f779d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[1]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[1]));
  AL_DFF_0 al_efd7be19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[2]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[2]));
  AL_DFF_0 al_ceb14878 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[11]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[11]));
  AL_DFF_0 al_d8a0a6b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[12]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[12]));
  AL_DFF_0 al_241e1370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[13]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[13]));
  AL_DFF_0 al_6969c7af (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[14]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[14]));
  AL_DFF_0 al_60758d0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[15]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[15]));
  AL_DFF_0 al_6079e76d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[16]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[16]));
  AL_DFF_0 al_9663f683 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[17]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[17]));
  AL_DFF_0 al_a7e566dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[44]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[44]));
  AL_DFF_0 al_5ed6db21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[45]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[45]));
  AL_DFF_0 al_b6590b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[46]),
    .en(al_a83e1130[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5c971b[46]));
  AL_DFF_0 al_9fb707a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[0]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[0]));
  AL_DFF_0 al_fead749 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[1]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[1]));
  AL_DFF_0 al_37e72e01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[2]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[2]));
  AL_DFF_0 al_10f150bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[11]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[11]));
  AL_DFF_0 al_70831f6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[12]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[12]));
  AL_DFF_0 al_9e0756da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[13]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[13]));
  AL_DFF_0 al_65c5313a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[14]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[14]));
  AL_DFF_0 al_9f0c2d89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[15]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[15]));
  AL_DFF_0 al_ef3b9b66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[16]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[16]));
  AL_DFF_0 al_4cea50c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[17]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[17]));
  AL_DFF_0 al_6a49e748 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[44]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[44]));
  AL_DFF_0 al_3e887e6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[45]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[45]));
  AL_DFF_0 al_6a686be9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8941a5fb[46]),
    .en(al_a83e1130[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51cc7f19[46]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    al_7392fa54 (
    .a(al_221aa358),
    .b(al_2dc3e45),
    .c(al_6ad3f77e),
    .d(al_369e229d[2]),
    .o(al_7c6fd728));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    al_62b3e7c4 (
    .a(al_7c6fd728),
    .b(al_8941a5fb[0]),
    .c(al_53bb123b[4]),
    .d(al_cbaa3056),
    .o(al_9bb5b978));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    al_a4a08cef (
    .a(al_7c6fd728),
    .b(al_8941a5fb[1]),
    .c(al_53bb123b[5]),
    .d(al_cbaa3056),
    .o(al_70777327));
  AL_DFF_0 al_725cfef7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9bb5b978),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53bb123b[4]));
  AL_DFF_0 al_b31fb165 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70777327),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53bb123b[5]));
  AL_DFF_0 al_b82b083b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e345b21[3]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_527755ec[3]));
  AL_DFF_0 al_7a30fd3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e345b21[4]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_527755ec[4]));
  AL_DFF_0 al_37ad76f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e345b21[0]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_527755ec[0]));
  AL_DFF_0 al_3423591e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e345b21[1]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_527755ec[1]));
  AL_DFF_0 al_9224fc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e345b21[2]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_527755ec[2]));
  AL_DFF_0 al_24b463d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[11]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2602b5cf[23]));
  AL_DFF_0 al_d0a647e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[12]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2602b5cf[24]));
  AL_DFF_0 al_9108b81c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[13]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2602b5cf[25]));
  AL_DFF_0 al_127279ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[14]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2602b5cf[26]));
  AL_DFF_0 al_95691798 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[15]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2602b5cf[27]));
  AL_DFF_0 al_cd0b03d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[16]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2602b5cf[28]));
  AL_DFF_0 al_e289ead9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e6e3a9da[17]),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_2602b5cf[29]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_cac90902 (
    .i(al_a3c26eaf),
    .o(al_82050a6e));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2679f086 (
    .i(al_82050a6e),
    .o(al_cbaa3056));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*B*~(C)*D*E)"),
    .INIT(32'h0800fbcf))
    al_4df497ef (
    .a(al_1d36bc6d),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_369e229d[2]),
    .e(al_7fb24d41[0]),
    .o(al_e048ecc8[0]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haacaa0aa))
    al_b5202581 (
    .a(al_e3f59f84[4]),
    .b(al_2a6634d6),
    .c(al_369e229d[0]),
    .d(al_369e229d[1]),
    .e(al_369e229d[2]),
    .o(al_e048ecc8[4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_55a27eca (
    .a(al_e048ecc8[4]),
    .b(al_e048ecc8[3]),
    .c(al_e048ecc8[2]),
    .d(al_e048ecc8[1]),
    .e(al_e048ecc8[0]),
    .o(al_1358d298));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~((F@E))+A*~(B)*~(C)*~(D)*~((F@E))+~(A)*B*~(C)*~(D)*~((F@E))+A*B*~(C)*~(D)*~((F@E))+~(A)*B*C*~(D)*~((F@E))+A*B*C*~(D)*~((F@E))+~(A)*~(B)*~(C)*D*~((F@E))+A*~(B)*~(C)*D*~((F@E))+A*B*~(C)*D*~((F@E))+~(A)*~(B)*C*D*~((F@E))+A*~(B)*C*D*~((F@E))+~(A)*B*C*D*~((F@E))+A*B*C*D*~((F@E))+A*B*~(C)*D*(F@E))"),
    .INIT(64'hfbcf08000800fbcf))
    al_87ad838c (
    .a(al_b0fb8887),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_369e229d[2]),
    .e(al_7fb24d41[0]),
    .f(al_7fb24d41[1]),
    .o(al_e048ecc8[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C@(~B*~A))"),
    .INIT(8'h1e))
    al_3ec3ea90 (
    .a(al_7fb24d41[0]),
    .b(al_7fb24d41[1]),
    .c(al_7fb24d41[2]),
    .o(al_8e600ada));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55c55055))
    al_e9ea6ad8 (
    .a(al_8e600ada),
    .b(al_a9552c76),
    .c(al_369e229d[0]),
    .d(al_369e229d[1]),
    .e(al_369e229d[2]),
    .o(al_e048ecc8[2]));
  AL_MAP_LUT4 #(
    .EQN("~(D@(~C*~B*~A))"),
    .INIT(16'h01fe))
    al_5876f830 (
    .a(al_7fb24d41[0]),
    .b(al_7fb24d41[1]),
    .c(al_7fb24d41[2]),
    .d(al_7fb24d41[3]),
    .o(al_629fa86a));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55c55055))
    al_4001547c (
    .a(al_629fa86a),
    .b(al_4331638),
    .c(al_369e229d[0]),
    .d(al_369e229d[1]),
    .e(al_369e229d[2]),
    .o(al_e048ecc8[3]));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~C*~B*~A))"),
    .INIT(32'hfffe0001))
    al_9c21048a (
    .a(al_7fb24d41[0]),
    .b(al_7fb24d41[1]),
    .c(al_7fb24d41[2]),
    .d(al_7fb24d41[3]),
    .e(al_7fb24d41[4]),
    .o(al_e3f59f84[4]));
  AL_DFF_0 al_9f30b56a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1358d298),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7e9a10b));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_80a303b3 (
    .a(al_9860067e),
    .b(al_f2dedfad[0]),
    .o(al_ca7553ae[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    al_b199f519 (
    .a(al_9860067e),
    .b(al_f2dedfad[0]),
    .c(al_f2dedfad[1]),
    .o(al_ca7553ae[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_e6a90cfd (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_ca7553ae[0]),
    .d(al_ca7553ae[1]),
    .o(al_3c502065));
  AL_DFF_0 al_c7b741c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3c502065),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9637b9));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b7d24d70 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[5]),
    .c(al_31adc4ab[0]),
    .o(al_10853ef5));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f3a1a1a3 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[5]),
    .c(al_39d4ac28[0]),
    .o(al_8c934a6b[0]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c485e1e3 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[5]),
    .c(al_2697e1b1[0]),
    .o(al_712e1022));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ede17991 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[5]),
    .c(al_f0541159[0]),
    .o(al_4084a330[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_8dfd2f31 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_10853ef5),
    .d(al_712e1022),
    .e(al_8c934a6b[0]),
    .f(al_4084a330[0]),
    .o(al_bc0d6480[0]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_5127da61 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[6]),
    .c(al_31adc4ab[11]),
    .o(al_9adb60d3));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_da7733f2 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[6]),
    .c(al_39d4ac28[11]),
    .o(al_8c934a6b[11]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e42d82cf (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[6]),
    .c(al_2697e1b1[11]),
    .o(al_a4dd1877));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_49709367 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[6]),
    .c(al_f0541159[11]),
    .o(al_4084a330[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_82c73b33 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_9adb60d3),
    .d(al_a4dd1877),
    .e(al_8c934a6b[11]),
    .f(al_4084a330[11]),
    .o(al_bc0d6480[11]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_66bb5c6a (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[7]),
    .c(al_31adc4ab[12]),
    .o(al_b7fe498b));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8702158b (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[7]),
    .c(al_39d4ac28[12]),
    .o(al_8c934a6b[12]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_539397c3 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[7]),
    .c(al_2697e1b1[12]),
    .o(al_d5de0442));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_912ac702 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[7]),
    .c(al_f0541159[12]),
    .o(al_4084a330[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_740a6678 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_b7fe498b),
    .d(al_d5de0442),
    .e(al_8c934a6b[12]),
    .f(al_4084a330[12]),
    .o(al_bc0d6480[12]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1ad4d8f (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[8]),
    .c(al_31adc4ab[13]),
    .o(al_b47d0925));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_eae74288 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[8]),
    .c(al_39d4ac28[13]),
    .o(al_8c934a6b[13]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_261806fd (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[8]),
    .c(al_2697e1b1[13]),
    .o(al_f4a06276));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_23a0c7fc (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[8]),
    .c(al_f0541159[13]),
    .o(al_4084a330[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_3c6cba8 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_b47d0925),
    .d(al_f4a06276),
    .e(al_8c934a6b[13]),
    .f(al_4084a330[13]),
    .o(al_bc0d6480[13]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c2ae2e4b (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[9]),
    .c(al_31adc4ab[14]),
    .o(al_a3e40416));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_93f6e5cb (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[9]),
    .c(al_39d4ac28[14]),
    .o(al_8c934a6b[14]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c42af17a (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[9]),
    .c(al_2697e1b1[14]),
    .o(al_8f975858));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_13f73e52 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[9]),
    .c(al_f0541159[14]),
    .o(al_4084a330[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_22e9b757 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_a3e40416),
    .d(al_8f975858),
    .e(al_8c934a6b[14]),
    .f(al_4084a330[14]),
    .o(al_bc0d6480[14]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_3bf2d394 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[10]),
    .c(al_31adc4ab[15]),
    .o(al_8b1b352d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_91ccc33a (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[10]),
    .c(al_39d4ac28[15]),
    .o(al_8c934a6b[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e0f88c3b (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[10]),
    .c(al_2697e1b1[15]),
    .o(al_7796e47d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_42a6e4b5 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[10]),
    .c(al_f0541159[15]),
    .o(al_4084a330[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_96a37845 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_8b1b352d),
    .d(al_7796e47d),
    .e(al_8c934a6b[15]),
    .f(al_4084a330[15]),
    .o(al_bc0d6480[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c5da0158 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[11]),
    .c(al_31adc4ab[16]),
    .o(al_a20b0983));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2228e22e (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[11]),
    .c(al_39d4ac28[16]),
    .o(al_8c934a6b[16]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_7a582cd6 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[11]),
    .c(al_2697e1b1[16]),
    .o(al_467e7732));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5020b637 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[11]),
    .c(al_f0541159[16]),
    .o(al_4084a330[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_33552a75 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_a20b0983),
    .d(al_467e7732),
    .e(al_8c934a6b[16]),
    .f(al_4084a330[16]),
    .o(al_bc0d6480[16]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b557ae67 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[12]),
    .c(al_31adc4ab[17]),
    .o(al_ea2829c1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_acc71fd6 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[12]),
    .c(al_39d4ac28[17]),
    .o(al_8c934a6b[17]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_68747acb (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[12]),
    .c(al_2697e1b1[17]),
    .o(al_e978fc5));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_65f24057 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[12]),
    .c(al_f0541159[17]),
    .o(al_4084a330[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_15840472 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_ea2829c1),
    .d(al_e978fc5),
    .e(al_8c934a6b[17]),
    .f(al_4084a330[17]),
    .o(al_bc0d6480[17]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_707a0937 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[3]),
    .c(al_2697e1b1[1]),
    .o(al_90f5a479));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_79dd1acf (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[3]),
    .c(al_f0541159[1]),
    .o(al_4084a330[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d1801dd4 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[3]),
    .c(al_39d4ac28[1]),
    .o(al_8c934a6b[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6dc3f93d (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[3]),
    .c(al_31adc4ab[1]),
    .o(al_6d99a7bb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haebf26378c9d0415))
    al_23b985dd (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_90f5a479),
    .d(al_6d99a7bb),
    .e(al_4084a330[1]),
    .f(al_8c934a6b[1]),
    .o(al_bc0d6480[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_7aa4c148 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[13]),
    .c(al_31adc4ab[24]),
    .o(al_37db4e3));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_41d13a33 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[13]),
    .c(al_39d4ac28[24]),
    .o(al_8c934a6b[24]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ddf0f54a (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[13]),
    .c(al_2697e1b1[24]),
    .o(al_4552d084));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_578f3b27 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[13]),
    .c(al_f0541159[24]),
    .o(al_4084a330[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_6b2d5deb (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_37db4e3),
    .d(al_4552d084),
    .e(al_8c934a6b[24]),
    .f(al_4084a330[24]),
    .o(al_bc0d6480[24]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1f624400 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[14]),
    .c(al_31adc4ab[25]),
    .o(al_be7cdff7));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e816ae7a (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[14]),
    .c(al_39d4ac28[25]),
    .o(al_8c934a6b[25]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ac7bd4e9 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[14]),
    .c(al_2697e1b1[25]),
    .o(al_50bc751d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d1df4191 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[14]),
    .c(al_f0541159[25]),
    .o(al_4084a330[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_9f114b54 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_be7cdff7),
    .d(al_50bc751d),
    .e(al_8c934a6b[25]),
    .f(al_4084a330[25]),
    .o(al_bc0d6480[25]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_730502aa (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[15]),
    .c(al_31adc4ab[26]),
    .o(al_374f7117));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_96a30455 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[15]),
    .c(al_39d4ac28[26]),
    .o(al_8c934a6b[26]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_539686d5 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[15]),
    .c(al_2697e1b1[26]),
    .o(al_169c4c39));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fdb59d01 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[15]),
    .c(al_f0541159[26]),
    .o(al_4084a330[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_a72bf224 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_374f7117),
    .d(al_169c4c39),
    .e(al_8c934a6b[26]),
    .f(al_4084a330[26]),
    .o(al_bc0d6480[26]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d6ff9f72 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[16]),
    .c(al_31adc4ab[27]),
    .o(al_ac0ca30d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_dd107add (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[16]),
    .c(al_39d4ac28[27]),
    .o(al_8c934a6b[27]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_626a5a53 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[16]),
    .c(al_2697e1b1[27]),
    .o(al_cec7db6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_cd5e3649 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[16]),
    .c(al_f0541159[27]),
    .o(al_4084a330[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_8aa03a9c (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_ac0ca30d),
    .d(al_cec7db6),
    .e(al_8c934a6b[27]),
    .f(al_4084a330[27]),
    .o(al_bc0d6480[27]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f9ca96d4 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[17]),
    .c(al_31adc4ab[28]),
    .o(al_7103149d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f15ad204 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[17]),
    .c(al_39d4ac28[28]),
    .o(al_8c934a6b[28]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_76012549 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[17]),
    .c(al_2697e1b1[28]),
    .o(al_b7ecdcb9));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d30ecaa4 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[17]),
    .c(al_f0541159[28]),
    .o(al_4084a330[28]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_e9641319 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_7103149d),
    .d(al_b7ecdcb9),
    .e(al_8c934a6b[28]),
    .f(al_4084a330[28]),
    .o(al_bc0d6480[28]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1f8913fe (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[18]),
    .c(al_31adc4ab[29]),
    .o(al_b55a64f2));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8f9c88e7 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[18]),
    .c(al_39d4ac28[29]),
    .o(al_8c934a6b[29]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9843f1b1 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[18]),
    .c(al_2697e1b1[29]),
    .o(al_95fc70f6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8492f543 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[18]),
    .c(al_f0541159[29]),
    .o(al_4084a330[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_7bce7361 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_b55a64f2),
    .d(al_95fc70f6),
    .e(al_8c934a6b[29]),
    .f(al_4084a330[29]),
    .o(al_bc0d6480[29]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b85633f4 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[4]),
    .c(al_31adc4ab[2]),
    .o(al_6f443675));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f1e9ce68 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[4]),
    .c(al_39d4ac28[2]),
    .o(al_8c934a6b[2]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b92bbd6d (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[4]),
    .c(al_2697e1b1[2]),
    .o(al_e72ab4a2));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1b20fb57 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[4]),
    .c(al_f0541159[2]),
    .o(al_4084a330[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_68e6ffb (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_6f443675),
    .d(al_e72ab4a2),
    .e(al_8c934a6b[2]),
    .f(al_4084a330[2]),
    .o(al_bc0d6480[2]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c4c3f628 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[19]),
    .c(al_31adc4ab[30]),
    .o(al_a6b23c82));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d15aeb2a (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[19]),
    .c(al_39d4ac28[30]),
    .o(al_8c934a6b[30]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a6926ef2 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[19]),
    .c(al_2697e1b1[30]),
    .o(al_51a643c1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3f1c667c (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[19]),
    .c(al_f0541159[30]),
    .o(al_4084a330[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_c76084be (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_a6b23c82),
    .d(al_51a643c1),
    .e(al_8c934a6b[30]),
    .f(al_4084a330[30]),
    .o(al_bc0d6480[30]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_8730d1aa (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[20]),
    .c(al_2697e1b1[31]),
    .o(al_4aab9ab7));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_504f24c6 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[20]),
    .c(al_f0541159[31]),
    .o(al_4084a330[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7c4fe92f (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[20]),
    .c(al_39d4ac28[31]),
    .o(al_8c934a6b[31]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_4895eb83 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[20]),
    .c(al_31adc4ab[31]),
    .o(al_2bdc9af8));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haebf26378c9d0415))
    al_2b3b1b4f (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_4aab9ab7),
    .d(al_2bdc9af8),
    .e(al_4084a330[31]),
    .f(al_8c934a6b[31]),
    .o(al_bc0d6480[31]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d2beab08 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[21]),
    .c(al_31adc4ab[32]),
    .o(al_5dbbae98));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3af475ee (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[21]),
    .c(al_39d4ac28[32]),
    .o(al_8c934a6b[32]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_878d7d66 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[21]),
    .c(al_2697e1b1[32]),
    .o(al_57c1f314));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_27ccab97 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[21]),
    .c(al_f0541159[32]),
    .o(al_4084a330[32]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_7f271f69 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_5dbbae98),
    .d(al_57c1f314),
    .e(al_8c934a6b[32]),
    .f(al_4084a330[32]),
    .o(al_bc0d6480[32]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_751185f8 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[22]),
    .c(al_31adc4ab[33]),
    .o(al_2aae8bdf));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_37d5a3c1 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[22]),
    .c(al_39d4ac28[33]),
    .o(al_8c934a6b[33]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1a490f80 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[22]),
    .c(al_2697e1b1[33]),
    .o(al_1370261a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bd3aedd5 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[22]),
    .c(al_f0541159[33]),
    .o(al_4084a330[33]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_884ae21d (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_2aae8bdf),
    .d(al_1370261a),
    .e(al_8c934a6b[33]),
    .f(al_4084a330[33]),
    .o(al_bc0d6480[33]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_468f855 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[23]),
    .c(al_31adc4ab[34]),
    .o(al_31640de4));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ab0ef64b (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[23]),
    .c(al_39d4ac28[34]),
    .o(al_8c934a6b[34]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_445aef88 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[23]),
    .c(al_2697e1b1[34]),
    .o(al_c3c25a23));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8e49a8dd (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[23]),
    .c(al_f0541159[34]),
    .o(al_4084a330[34]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_d835de1c (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_31640de4),
    .d(al_c3c25a23),
    .e(al_8c934a6b[34]),
    .f(al_4084a330[34]),
    .o(al_bc0d6480[34]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_817276d9 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[24]),
    .c(al_31adc4ab[35]),
    .o(al_e5b96d96));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e958451c (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[24]),
    .c(al_39d4ac28[35]),
    .o(al_8c934a6b[35]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ceb19bf7 (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[24]),
    .c(al_2697e1b1[35]),
    .o(al_bd7030bd));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_dff8aaf5 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[24]),
    .c(al_f0541159[35]),
    .o(al_4084a330[35]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_32f7a020 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_e5b96d96),
    .d(al_bd7030bd),
    .e(al_8c934a6b[35]),
    .f(al_4084a330[35]),
    .o(al_bc0d6480[35]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_fe5d03c7 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[25]),
    .c(al_31adc4ab[36]),
    .o(al_69e722f9));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4d57d640 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[25]),
    .c(al_39d4ac28[36]),
    .o(al_8c934a6b[36]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f1ef39fb (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[25]),
    .c(al_2697e1b1[36]),
    .o(al_7f1ab5ea));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_faa102d7 (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[25]),
    .c(al_f0541159[36]),
    .o(al_4084a330[36]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_b99087ed (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_69e722f9),
    .d(al_7f1ab5ea),
    .e(al_8c934a6b[36]),
    .f(al_4084a330[36]),
    .o(al_bc0d6480[36]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c8f3124 (
    .a(al_ef92c438[0]),
    .b(al_58fb4752[26]),
    .c(al_31adc4ab[37]),
    .o(al_2f16accf));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_69670bc5 (
    .a(al_ef92c438[1]),
    .b(al_58fb4752[26]),
    .c(al_39d4ac28[37]),
    .o(al_8c934a6b[37]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_446e4b6f (
    .a(al_ef92c438[2]),
    .b(al_58fb4752[26]),
    .c(al_2697e1b1[37]),
    .o(al_1dbbf5ed));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7d76c3ae (
    .a(al_ef92c438[3]),
    .b(al_58fb4752[26]),
    .c(al_f0541159[37]),
    .o(al_4084a330[37]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_d3200ca9 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_2f16accf),
    .d(al_1dbbf5ed),
    .e(al_8c934a6b[37]),
    .f(al_4084a330[37]),
    .o(al_bc0d6480[37]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_cef2bf74 (
    .a(al_ef92c438[0]),
    .b(al_88a8db2c[0]),
    .c(al_31adc4ab[44]),
    .o(al_6e1be86c));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_250c203a (
    .a(al_ef92c438[1]),
    .b(al_88a8db2c[0]),
    .c(al_39d4ac28[44]),
    .o(al_8c934a6b[44]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_2d7b151c (
    .a(al_ef92c438[2]),
    .b(al_88a8db2c[0]),
    .c(al_2697e1b1[44]),
    .o(al_3a4ffd2d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_61577dd5 (
    .a(al_ef92c438[3]),
    .b(al_88a8db2c[0]),
    .c(al_f0541159[44]),
    .o(al_4084a330[44]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_67f8eab2 (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_6e1be86c),
    .d(al_3a4ffd2d),
    .e(al_8c934a6b[44]),
    .f(al_4084a330[44]),
    .o(al_bc0d6480[44]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a773b75e (
    .a(al_ef92c438[0]),
    .b(al_88a8db2c[1]),
    .c(al_31adc4ab[45]),
    .o(al_ac21ff42));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f5645e00 (
    .a(al_ef92c438[1]),
    .b(al_88a8db2c[1]),
    .c(al_39d4ac28[45]),
    .o(al_8c934a6b[45]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f53db6ab (
    .a(al_ef92c438[2]),
    .b(al_88a8db2c[1]),
    .c(al_2697e1b1[45]),
    .o(al_5e53d63d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_432f91bd (
    .a(al_ef92c438[3]),
    .b(al_88a8db2c[1]),
    .c(al_f0541159[45]),
    .o(al_4084a330[45]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_be4aad3c (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_ac21ff42),
    .d(al_5e53d63d),
    .e(al_8c934a6b[45]),
    .f(al_4084a330[45]),
    .o(al_bc0d6480[45]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_38c2686f (
    .a(al_ca7553ae[0]),
    .b(al_f2dedfad[1]),
    .o(al_ef92c438[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c68f525a (
    .a(al_ef92c438[3]),
    .b(al_88a8db2c[2]),
    .c(al_f0541159[46]),
    .o(al_4084a330[46]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_a24dc2ed (
    .a(al_b528368c[0]),
    .b(al_b528368c[1]),
    .c(al_70c05302),
    .d(al_392853fb),
    .e(al_8c934a6b[46]),
    .f(al_4084a330[46]),
    .o(al_bc0d6480[46]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_405ee49f (
    .a(al_ca7553ae[0]),
    .b(al_ca7553ae[1]),
    .o(al_ef92c438[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_c7b768b6 (
    .a(al_ca7553ae[0]),
    .b(al_ca7553ae[1]),
    .o(al_ef92c438[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5a15a639 (
    .a(al_ca7553ae[0]),
    .b(al_f2dedfad[1]),
    .o(al_ef92c438[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_9887e7c6 (
    .a(al_ef92c438[0]),
    .b(al_88a8db2c[2]),
    .c(al_31adc4ab[46]),
    .o(al_70c05302));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_982fcce6 (
    .a(al_ef92c438[1]),
    .b(al_88a8db2c[2]),
    .c(al_39d4ac28[46]),
    .o(al_8c934a6b[46]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1947c37c (
    .a(al_ef92c438[2]),
    .b(al_88a8db2c[2]),
    .c(al_2697e1b1[46]),
    .o(al_392853fb));
  AL_DFF_0 al_3fc63ded (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55876a5e),
    .en(1'b1),
    .sr(al_cbaa3056),
    .ss(1'b0),
    .q(al_f419b7f2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_b65aa411 (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[0]),
    .d(al_e9ebbe15[0]),
    .e(al_c5c971b[0]),
    .f(al_51cc7f19[0]),
    .o(al_9b520651));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_e18303c5 (
    .a(al_369e229d[0]),
    .b(al_369e229d[1]),
    .o(al_6ad3f77e));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_88d3bc75 (
    .a(al_403fbf52),
    .b(al_53439d34),
    .c(al_8941a5fb[0]),
    .o(al_524a1bfd));
  AL_MAP_LUT6 #(
    .EQN("(F@~(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'hf0cc55550f33aaaa))
    al_fea74e6d (
    .a(al_524a1bfd),
    .b(al_2a5fa8c),
    .c(al_ebe69372),
    .d(al_8941a5fb[0]),
    .e(al_8941a5fb[1]),
    .f(al_8941a5fb[35]),
    .o(al_dfc3cb3c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_93f1d3d1 (
    .a(al_a4914504),
    .b(al_a1d2ac98),
    .c(al_34ff0ff5),
    .d(al_18d4d578),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_87136fec));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_48026885 (
    .a(al_3185ed47),
    .b(al_bfe0071c),
    .c(al_6692b66c),
    .d(al_e80539a7),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_416ad84c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_c72ee81d (
    .a(al_e2bcb10),
    .b(al_25de7719),
    .c(al_49d43cfa),
    .d(al_fc1936a5),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_cb0fcfc7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_b52d2c8b (
    .a(al_b1edca88),
    .b(al_364b2d93),
    .c(al_28da8a0d),
    .d(al_e1521e17),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_b2365485));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_74042c2a (
    .a(al_2e96480),
    .b(al_22a3e261),
    .c(al_3647cd0),
    .d(al_9526df3b),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_7eb31edc));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_fc7e17cc (
    .a(al_9d701591),
    .b(al_bd5f3c97),
    .c(al_e4c2295a),
    .d(al_26b95353),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_bdded574));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_425b10b4 (
    .a(al_9264d6ce),
    .b(al_9dee74a8),
    .c(al_8941a5fb[0]),
    .o(al_8a3c47e1));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_67eda969 (
    .a(al_9b520651),
    .b(al_9e2903f5),
    .c(al_8941a5fb[0]),
    .o(al_e6e3a9da[0]));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_623e623f (
    .a(al_8a3c47e1),
    .b(al_b62c6ace),
    .c(al_c959a932),
    .d(al_8941a5fb[0]),
    .e(al_8941a5fb[1]),
    .f(al_8941a5fb[31]),
    .o(al_631e0c37));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_cc25fd72 (
    .a(al_48aee091),
    .b(al_10d1f7da),
    .c(al_539c7732),
    .d(al_a448873e),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_3a3118b0));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_689fb59 (
    .a(al_1b6a0af9),
    .b(al_6a2ba50d),
    .c(al_8941a5fb[0]),
    .o(al_d8ecb3f8));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_d3036d9f (
    .a(al_d8ecb3f8),
    .b(al_c32d8f29),
    .c(al_66bed231),
    .d(al_8941a5fb[0]),
    .e(al_8941a5fb[1]),
    .f(al_8941a5fb[33]),
    .o(al_bd4dc0cb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_e3fa7ac5 (
    .a(al_464fb058),
    .b(al_fd5ac0c0),
    .c(al_6bbd7053),
    .d(al_dd9df6a3),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_d6e5ffe2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_56adcf58 (
    .a(al_e707cc02),
    .b(al_e2740cd5),
    .c(al_4743871),
    .d(al_f498aaed),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_c092a1dc));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_dd40b039 (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[1]),
    .d(al_e9ebbe15[1]),
    .e(al_c5c971b[1]),
    .f(al_51cc7f19[1]),
    .o(al_9c060979));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_69429802 (
    .a(al_5d3dfa86),
    .b(al_55c1f3f8),
    .c(al_2f5e01b7),
    .d(al_a04a63d4),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_995c4dc4));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_9dfb5a62 (
    .a(al_8287cea7),
    .b(al_dedd5989),
    .c(al_8941a5fb[0]),
    .o(al_b7abf9db));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_bc906544 (
    .a(al_b7abf9db),
    .b(al_b4d9e182),
    .c(al_e0a71537),
    .d(al_8941a5fb[0]),
    .e(al_8941a5fb[1]),
    .f(al_8941a5fb[36]),
    .o(al_846eafad));
  AL_MAP_LUT6 #(
    .EQN("((D@C)*(F@B)*(E@A))"),
    .INIT(64'h0110022004400880))
    al_ed451157 (
    .a(al_bdded574),
    .b(al_3a3118b0),
    .c(al_c092a1dc),
    .d(al_8941a5fb[24]),
    .e(al_8941a5fb[26]),
    .f(al_8941a5fb[28]),
    .o(al_7b43c1e));
  AL_MAP_LUT6 #(
    .EQN("(~B*A*(E@D)*(F@C))"),
    .INIT(64'h0002020000202000))
    al_c719bcde (
    .a(al_dfc3cb3c),
    .b(al_846eafad),
    .c(al_cb0fcfc7),
    .d(al_7eb31edc),
    .e(al_8941a5fb[30]),
    .f(al_8941a5fb[32]),
    .o(al_6860fc86));
  AL_MAP_LUT6 #(
    .EQN("((D@C)*(E@B)*(F@A))"),
    .INIT(64'h0110044002200880))
    al_6411f6 (
    .a(al_416ad84c),
    .b(al_b2365485),
    .c(al_d6e5ffe2),
    .d(al_8941a5fb[25]),
    .e(al_8941a5fb[27]),
    .f(al_8941a5fb[29]),
    .o(al_8cddf958));
  AL_MAP_LUT6 #(
    .EQN("(~B*~A*(E@D)*(F@C))"),
    .INIT(64'h0001010000101000))
    al_e722201e (
    .a(al_631e0c37),
    .b(al_bd4dc0cb),
    .c(al_87136fec),
    .d(al_995c4dc4),
    .e(al_8941a5fb[34]),
    .f(al_8941a5fb[37]),
    .o(al_74055ffa));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_e2d6e147 (
    .a(al_833f5c05),
    .b(al_3df83ccd),
    .c(al_61792012),
    .d(al_286587c2),
    .e(al_8941a5fb[0]),
    .f(al_8941a5fb[1]),
    .o(al_c711503f));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*~B))"),
    .INIT(16'h0405))
    al_27a8fa10 (
    .a(al_c711503f),
    .b(al_9860067e),
    .c(al_79dddfae),
    .d(al_ad9637b9),
    .o(al_f027c275));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_f185dcd9 (
    .a(al_6860fc86),
    .b(al_74055ffa),
    .c(al_7b43c1e),
    .d(al_8cddf958),
    .e(al_f027c275),
    .f(al_6ad3f77e),
    .o(al_cefb896));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(E*C*B*~A))"),
    .INIT(32'h00bf00ff))
    al_c0633a64 (
    .a(al_79dddfae),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_369e229d[2]),
    .e(al_c360bf4c[2]),
    .o(al_485702b6));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_267b807 (
    .a(al_9c060979),
    .b(al_9e2903f5),
    .c(al_8941a5fb[1]),
    .o(al_e6e3a9da[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_36b1a923 (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[45]),
    .d(al_e9ebbe15[45]),
    .e(al_c5c971b[45]),
    .f(al_51cc7f19[45]),
    .o(al_fa2c6203));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_68627b95 (
    .a(al_fa2c6203),
    .b(al_9e2903f5),
    .c(al_8941a5fb[45]),
    .o(al_e6a713a5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_e664cc6a (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[46]),
    .d(al_e9ebbe15[46]),
    .e(al_c5c971b[46]),
    .f(al_51cc7f19[46]),
    .o(al_2d84af31));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_aece4e2e (
    .a(al_2d84af31),
    .b(al_9e2903f5),
    .c(al_8941a5fb[46]),
    .o(al_e6e3a9da[46]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_3d952062 (
    .a(al_11a7c870[0]),
    .b(al_11a7c870[1]),
    .c(al_59b0cd05[44]),
    .d(al_e9ebbe15[44]),
    .e(al_c5c971b[44]),
    .f(al_51cc7f19[44]),
    .o(al_a807c60d));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_f7ecbbc2 (
    .a(al_a807c60d),
    .b(al_9e2903f5),
    .c(al_8941a5fb[44]),
    .o(al_3e892816));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_60400d98 (
    .a(init_calib_complete),
    .b(al_90d84dc7[2]),
    .c(al_61f44420),
    .d(ddr_app_rdy),
    .o(al_9860067e));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_64ca5d09 (
    .a(al_e6e3a9da[46]),
    .b(al_3e892816),
    .o(al_732fadca));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_37cda037 (
    .a(al_e6e3a9da[0]),
    .b(al_e6e3a9da[1]),
    .c(al_1cf815c1),
    .d(al_c74d7793),
    .e(al_82bb1e86),
    .f(al_3b347f86),
    .o(al_84bf2198));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~(~D*~(C*~A))))"),
    .INIT(32'h00233333))
    al_86df1fc0 (
    .a(al_cefb896),
    .b(al_84bf2198),
    .c(al_485702b6),
    .d(al_13f9c71c),
    .e(al_9e2903f5),
    .o(al_85567015));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_d9a22c0 (
    .a(al_732fadca),
    .b(al_e6a713a5),
    .o(al_b3701730));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_484aa85 (
    .a(al_e6a713a5),
    .b(al_e6e3a9da[46]),
    .c(al_3e892816),
    .d(al_1f97cafb[0]),
    .e(al_1f97cafb[1]),
    .o(al_f748e656));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~(C*~B*A)))"),
    .INIT(32'h00ff0020))
    al_1b09444e (
    .a(al_85567015),
    .b(al_b3701730),
    .c(al_f748e656),
    .d(al_ef78cbcb),
    .e(al_f419b7f2),
    .o(al_55876a5e));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    al_bf9c3f09 (
    .a(al_79dddfae),
    .b(al_369e229d[0]),
    .c(al_369e229d[1]),
    .d(al_369e229d[2]),
    .o(al_13f9c71c));
  AL_DFF_0 al_a95b995e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c4726cab),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90d84dc7[3]));
  AL_DFF_0 al_de215051 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f4cc2ce5),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_1c8747c7));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e2c3a8dc (
    .a(al_3e56391),
    .b(al_12521532),
    .o(al_321810b0));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_bbc06ad2 (
    .a(al_465b8d7d),
    .b(al_c360bf4c[3]),
    .o(al_f4cc2ce5));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_f43ec236 (
    .a(al_ef35f7b6[0]),
    .b(al_ef35f7b6[1]),
    .c(al_b25d0e99[1]),
    .d(al_fea7bbd9[0]),
    .e(al_fea7bbd9[1]),
    .o(al_9941ff24[1]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_ae6e78ae (
    .a(al_ef35f7b6[0]),
    .b(al_ef35f7b6[1]),
    .c(al_b25d0e99[2]),
    .d(al_16b7523e[0]),
    .e(al_16b7523e[1]),
    .o(al_9941ff24[2]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E@B)*~(D@A))"),
    .INIT(32'h80402010))
    al_108a2b2c (
    .a(al_ef35f7b6[0]),
    .b(al_ef35f7b6[1]),
    .c(al_b25d0e99[0]),
    .d(al_974136cc[0]),
    .e(al_974136cc[1]),
    .o(al_9941ff24[0]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(D*~(F@C)*~(E@B)))"),
    .INIT(64'h1555455551555455))
    al_fec670ef (
    .a(al_9941ff24[2]),
    .b(al_ef35f7b6[0]),
    .c(al_ef35f7b6[1]),
    .d(al_b25d0e99[3]),
    .e(al_f82ace94[0]),
    .f(al_f82ace94[1]),
    .o(al_65e4d4e0));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_70f7183f (
    .a(al_65e4d4e0),
    .b(al_321810b0),
    .c(al_82001be8),
    .d(al_9941ff24[1]),
    .e(al_9941ff24[0]),
    .o(al_65bd6ac6));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(~D*(A*C*~(E)*~(F)+A*C*~(E)*F+~(A)*~(C)*E*F+A*~(C)*E*F)))"),
    .INIT(64'h3330331333333313))
    al_9939ede9 (
    .a(al_65bd6ac6),
    .b(al_1c8747c7),
    .c(al_9d2be50d[0]),
    .d(al_9d2be50d[1]),
    .e(al_9d2be50d[2]),
    .f(al_530cb84f),
    .o(al_465b8d7d));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*~A))"),
    .INIT(8'hc9))
    al_9009c54c (
    .a(al_1a411806),
    .b(al_6ea52063),
    .c(al_c28589ac),
    .o(al_f6114766[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(~D*~B*~A))"),
    .INIT(16'hf0e1))
    al_8db7187c (
    .a(al_1a411806),
    .b(al_6ea52063),
    .c(al_4d29fbf3),
    .d(al_c28589ac),
    .o(al_f6114766[2]));
  AL_MAP_LUT6 #(
    .EQN("(E@(~F*~D*~C*~B*~A))"),
    .INIT(64'hffff0000fffe0001))
    al_1ee6c7c6 (
    .a(al_1a411806),
    .b(al_6ea52063),
    .c(al_4d29fbf3),
    .d(al_f2c5bff2),
    .e(al_862761d2),
    .f(al_c28589ac),
    .o(al_f6114766[4]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_ee7ab428 (
    .a(al_1a411806),
    .b(al_c28589ac),
    .o(al_f6114766[0]));
  AL_MAP_LUT5 #(
    .EQN("(D@(~E*~C*~B*~A))"),
    .INIT(32'hff00fe01))
    al_2a5decc7 (
    .a(al_1a411806),
    .b(al_6ea52063),
    .c(al_4d29fbf3),
    .d(al_f2c5bff2),
    .e(al_c28589ac),
    .o(al_f6114766[3]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_e2268020 (
    .a(al_f6114766[3]),
    .b(al_f6114766[0]),
    .c(al_6ea52063),
    .d(al_4d29fbf3),
    .e(al_862761d2),
    .o(al_9c4fa309[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_a4a2ce5e (
    .a(al_9c4fa309[0]),
    .b(al_c28589ac),
    .o(al_71faa803[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_39825b7d (
    .a(al_dd768853[0]),
    .b(al_eec54698[0]),
    .c(al_ffdc699f[0]),
    .d(al_f1974c03[0]),
    .e(al_a196b5f4[0]),
    .f(al_a196b5f4[1]),
    .o(al_a3f7dedc[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_f1e1c83e (
    .a(al_dd768853[1]),
    .b(al_eec54698[1]),
    .c(al_ffdc699f[1]),
    .d(al_f1974c03[1]),
    .e(al_a196b5f4[0]),
    .f(al_a196b5f4[1]),
    .o(al_a3f7dedc[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_1a39e17b (
    .a(al_dd768853[2]),
    .b(al_eec54698[2]),
    .c(al_ffdc699f[2]),
    .d(al_f1974c03[2]),
    .e(al_a196b5f4[0]),
    .f(al_a196b5f4[1]),
    .o(al_a3f7dedc[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_f65d87 (
    .a(al_dd768853[3]),
    .b(al_eec54698[3]),
    .c(al_ffdc699f[3]),
    .d(al_f1974c03[3]),
    .e(al_a196b5f4[0]),
    .f(al_a196b5f4[1]),
    .o(al_a3f7dedc[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_497ca040 (
    .a(al_dd768853[4]),
    .b(al_eec54698[4]),
    .c(al_ffdc699f[4]),
    .d(al_f1974c03[4]),
    .e(al_a196b5f4[0]),
    .f(al_a196b5f4[1]),
    .o(al_a3f7dedc[4]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    al_b0dfd (
    .a(al_d51c2ed1),
    .b(al_10aff3dd[0]),
    .c(al_10aff3dd[1]),
    .o(al_b97c37dd));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_13669183 (
    .a(al_b97c37dd),
    .b(al_a196b5f4[0]),
    .o(al_68f1a7a7[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*~A))"),
    .INIT(8'hb4))
    al_20ae6256 (
    .a(al_b97c37dd),
    .b(al_a196b5f4[0]),
    .c(al_a196b5f4[1]),
    .o(al_68f1a7a7[1]));
  AL_MAP_LUT4 #(
    .EQN("(D@(~C*~(B*~A)))"),
    .INIT(16'hf40b))
    al_e6fcb27f (
    .a(al_d7badb25),
    .b(al_c693d245),
    .c(al_edebd92e),
    .d(al_b1a73cf[0]),
    .o(al_e11b20ed[0]));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~C*~(B*~A)))"),
    .INIT(32'hf4ff0b00))
    al_426a0d79 (
    .a(al_d7badb25),
    .b(al_c693d245),
    .c(al_edebd92e),
    .d(al_b1a73cf[0]),
    .e(al_b1a73cf[1]),
    .o(al_e11b20ed[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_3a928dcd (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_68f1a7a7[0]),
    .d(al_68f1a7a7[1]),
    .o(al_21409483));
  AL_DFF_0 al_bcbbedb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21409483),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d149d704));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(C*~A))"),
    .INIT(16'h639c))
    al_df37db3b (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_68f1a7a7[0]),
    .d(al_68f1a7a7[1]),
    .o(al_eacb80c[1]));
  AL_DFF_0 al_6048dc7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eacb80c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c088e9dc));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_922b8b1b (
    .a(al_b1a73cf[0]),
    .b(al_b1a73cf[1]),
    .o(al_69c2ff54[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(~E*~D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffffffcca0a0a080))
    al_e6c8bd97 (
    .a(al_ec7a421c),
    .b(al_b97c37dd),
    .c(al_69c2ff54[0]),
    .d(al_a196b5f4[0]),
    .e(al_a196b5f4[1]),
    .f(al_b25d0e99[0]),
    .o(al_696c7934[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5caed2e6 (
    .a(al_b1a73cf[0]),
    .b(al_b1a73cf[1]),
    .o(al_69c2ff54[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(~E*D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffffccffa0a080a0))
    al_eb67f71f (
    .a(al_ec7a421c),
    .b(al_b97c37dd),
    .c(al_69c2ff54[1]),
    .d(al_a196b5f4[0]),
    .e(al_a196b5f4[1]),
    .f(al_b25d0e99[1]),
    .o(al_696c7934[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_da6509d1 (
    .a(al_b1a73cf[0]),
    .b(al_b1a73cf[1]),
    .o(al_69c2ff54[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(E*~D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hffccffffa080a0a0))
    al_32354d34 (
    .a(al_ec7a421c),
    .b(al_b97c37dd),
    .c(al_69c2ff54[2]),
    .d(al_a196b5f4[0]),
    .e(al_a196b5f4[1]),
    .f(al_b25d0e99[2]),
    .o(al_696c7934[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_6e57b2ff (
    .a(al_b1a73cf[0]),
    .b(al_b1a73cf[1]),
    .o(al_69c2ff54[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    al_939b3970 (
    .a(al_d7badb25),
    .b(al_c693d245),
    .c(al_edebd92e),
    .o(al_ec7a421c));
  AL_MAP_LUT6 #(
    .EQN("(~(E*D*~B)*~(~F*~(C*A)))"),
    .INIT(64'hccffffff80a0a0a0))
    al_d3bbd5d1 (
    .a(al_ec7a421c),
    .b(al_b97c37dd),
    .c(al_69c2ff54[3]),
    .d(al_a196b5f4[0]),
    .e(al_a196b5f4[1]),
    .f(al_b25d0e99[3]),
    .o(al_696c7934[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_35a86c5e (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[11]),
    .d(al_fea7bbd9[11]),
    .e(al_16b7523e[11]),
    .f(al_f82ace94[11]),
    .o(al_4a34f384));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_709fa1c0 (
    .a(al_4a34f384),
    .b(al_d149d704),
    .c(al_ef35f7b6[11]),
    .o(al_7040e81f[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_74d56a87 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[12]),
    .d(al_fea7bbd9[12]),
    .e(al_16b7523e[12]),
    .f(al_f82ace94[12]),
    .o(al_90420b48));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_df52e3ba (
    .a(al_90420b48),
    .b(al_d149d704),
    .c(al_ef35f7b6[12]),
    .o(al_7040e81f[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_734f1d23 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[13]),
    .d(al_fea7bbd9[13]),
    .e(al_16b7523e[13]),
    .f(al_f82ace94[13]),
    .o(al_3f896a8c));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_6841f7ce (
    .a(al_3f896a8c),
    .b(al_d149d704),
    .c(al_ef35f7b6[13]),
    .o(al_7040e81f[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_b3fb4388 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[14]),
    .d(al_fea7bbd9[14]),
    .e(al_16b7523e[14]),
    .f(al_f82ace94[14]),
    .o(al_177ed223));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_6f27c8c2 (
    .a(al_177ed223),
    .b(al_d149d704),
    .c(al_ef35f7b6[14]),
    .o(al_7040e81f[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_2a2b4f3f (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[15]),
    .d(al_fea7bbd9[15]),
    .e(al_16b7523e[15]),
    .f(al_f82ace94[15]),
    .o(al_af2a474d));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_2aad1423 (
    .a(al_af2a474d),
    .b(al_d149d704),
    .c(al_ef35f7b6[15]),
    .o(al_7040e81f[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_219675aa (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[16]),
    .d(al_fea7bbd9[16]),
    .e(al_16b7523e[16]),
    .f(al_f82ace94[16]),
    .o(al_8dcb6b40));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_3a16fa3b (
    .a(al_8dcb6b40),
    .b(al_d149d704),
    .c(al_ef35f7b6[16]),
    .o(al_7040e81f[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_2b3f2d81 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[17]),
    .d(al_fea7bbd9[17]),
    .e(al_16b7523e[17]),
    .f(al_f82ace94[17]),
    .o(al_5b157bf));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_37a907dd (
    .a(al_5b157bf),
    .b(al_d149d704),
    .c(al_ef35f7b6[17]),
    .o(al_7040e81f[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_9b98fe45 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[2]),
    .d(al_fea7bbd9[2]),
    .e(al_16b7523e[2]),
    .f(al_f82ace94[2]),
    .o(al_a4747624));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_67b3cae0 (
    .a(al_a4747624),
    .b(al_d149d704),
    .c(al_ef35f7b6[2]),
    .o(al_7040e81f[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_bb1c7db3 (
    .a(al_89ad3a7d[0]),
    .b(al_45d9e18e[0]),
    .c(al_c5e4c82d[0]),
    .d(al_9892447e[0]),
    .e(al_1124d2df[0]),
    .f(al_1124d2df[1]),
    .o(al_bf99db4a));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_bdb26f59 (
    .a(al_bf99db4a),
    .b(al_3e56391),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[0]),
    .f(al_75c0d27f[0]),
    .o(al_b671fee2[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_20f5b17 (
    .a(al_b671fee2[0]),
    .b(al_45d9e18e[0]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_c325b022[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_452203bd (
    .a(al_b671fee2[0]),
    .b(al_9892447e[0]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_1a25e1aa[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_d88a8b3c (
    .a(al_b671fee2[0]),
    .b(al_c5e4c82d[0]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_6f7a76fc[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_a888b456 (
    .a(al_b671fee2[0]),
    .b(al_89ad3a7d[0]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_2497ff95[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_76de918b (
    .a(al_c325b022[0]),
    .b(al_1a25e1aa[0]),
    .c(al_6f7a76fc[0]),
    .d(al_2497ff95[0]),
    .e(al_b1a73cf[0]),
    .f(al_b1a73cf[1]),
    .o(al_5b784e0e[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_f4c200e (
    .a(al_89ad3a7d[1]),
    .b(al_45d9e18e[1]),
    .c(al_c5e4c82d[1]),
    .d(al_9892447e[1]),
    .e(al_1124d2df[0]),
    .f(al_1124d2df[1]),
    .o(al_e76a8396));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'h22222ee2e22eeeee))
    al_18bbd24e (
    .a(al_e76a8396),
    .b(al_3e56391),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[1]),
    .f(al_75c0d27f[1]),
    .o(al_e5a22863));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((~D*C))+~B*A*~((~D*C))+~(~B)*A*(~D*C)+~B*A*(~D*C))"),
    .INIT(16'hcc5c))
    al_336678d1 (
    .a(al_e5a22863),
    .b(al_45d9e18e[1]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_c325b022[1]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((D*C))+~B*A*~((D*C))+~(~B)*A*(D*C)+~B*A*(D*C))"),
    .INIT(16'h5ccc))
    al_d61f82c (
    .a(al_e5a22863),
    .b(al_9892447e[1]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_1a25e1aa[1]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((D*~C))+~B*A*~((D*~C))+~(~B)*A*(D*~C)+~B*A*(D*~C))"),
    .INIT(16'hc5cc))
    al_24abf197 (
    .a(al_e5a22863),
    .b(al_c5e4c82d[1]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_6f7a76fc[1]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A)*~((~D*~C))+~B*A*~((~D*~C))+~(~B)*A*(~D*~C)+~B*A*(~D*~C))"),
    .INIT(16'hccc5))
    al_8afc92a8 (
    .a(al_e5a22863),
    .b(al_89ad3a7d[1]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_2497ff95[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_8fcfb539 (
    .a(al_c325b022[1]),
    .b(al_1a25e1aa[1]),
    .c(al_6f7a76fc[1]),
    .d(al_2497ff95[1]),
    .e(al_b1a73cf[0]),
    .f(al_b1a73cf[1]),
    .o(al_5b784e0e[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_4d44b1c8 (
    .a(al_89ad3a7d[2]),
    .b(al_45d9e18e[2]),
    .c(al_c5e4c82d[2]),
    .d(al_9892447e[2]),
    .e(al_1124d2df[0]),
    .f(al_1124d2df[1]),
    .o(al_39f329dd));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_d2309415 (
    .a(al_39f329dd),
    .b(al_3e56391),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[2]),
    .f(al_75c0d27f[2]),
    .o(al_b671fee2[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_a2cb2feb (
    .a(al_b671fee2[2]),
    .b(al_45d9e18e[2]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_c325b022[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_3b023122 (
    .a(al_b671fee2[2]),
    .b(al_9892447e[2]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_1a25e1aa[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_62ed6eb9 (
    .a(al_b671fee2[2]),
    .b(al_c5e4c82d[2]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_6f7a76fc[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_6af40874 (
    .a(al_b671fee2[2]),
    .b(al_89ad3a7d[2]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_2497ff95[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_6b9ea6cb (
    .a(al_c325b022[2]),
    .b(al_1a25e1aa[2]),
    .c(al_6f7a76fc[2]),
    .d(al_2497ff95[2]),
    .e(al_b1a73cf[0]),
    .f(al_b1a73cf[1]),
    .o(al_5b784e0e[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_34b0934c (
    .a(al_89ad3a7d[3]),
    .b(al_45d9e18e[3]),
    .c(al_c5e4c82d[3]),
    .d(al_9892447e[3]),
    .e(al_1124d2df[0]),
    .f(al_1124d2df[1]),
    .o(al_73c5a4c));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C)))*~(B)+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*~(B)+~(~A)*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B+~A*(F*~(E)*~((D@C))+F*E*~((D@C))+~(F)*E*(D@C)+F*E*(D@C))*B)"),
    .INIT(64'hddddd11d1dd11111))
    al_21dcdf69 (
    .a(al_73c5a4c),
    .b(al_3e56391),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[3]),
    .f(al_75c0d27f[3]),
    .o(al_b671fee2[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_3c79f18c (
    .a(al_b671fee2[3]),
    .b(al_45d9e18e[3]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_c325b022[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_79c408af (
    .a(al_b671fee2[3]),
    .b(al_9892447e[3]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_1a25e1aa[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_409ed37e (
    .a(al_b671fee2[3]),
    .b(al_c5e4c82d[3]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_6f7a76fc[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_6b2c7610 (
    .a(al_b671fee2[3]),
    .b(al_89ad3a7d[3]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_2497ff95[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_845712eb (
    .a(al_c325b022[3]),
    .b(al_1a25e1aa[3]),
    .c(al_6f7a76fc[3]),
    .d(al_2497ff95[3]),
    .e(al_b1a73cf[0]),
    .f(al_b1a73cf[1]),
    .o(al_5b784e0e[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_34152442 (
    .a(al_89ad3a7d[4]),
    .b(al_45d9e18e[4]),
    .c(al_c5e4c82d[4]),
    .d(al_9892447e[4]),
    .e(al_1124d2df[0]),
    .f(al_1124d2df[1]),
    .o(al_60eb3a40));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*(D@C)))*~(B)+~A*(E*(D@C))*~(B)+~(~A)*(E*(D@C))*B+~A*(E*(D@C))*B)"),
    .INIT(32'h1dd11111))
    al_677502ad (
    .a(al_60eb3a40),
    .b(al_3e56391),
    .c(al_bfd664bf[0]),
    .d(al_bfd664bf[1]),
    .e(al_17e51133[4]),
    .o(al_b671fee2[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*C))+B*A*~((~D*C))+~(B)*A*(~D*C)+B*A*(~D*C))"),
    .INIT(16'hccac))
    al_9d809050 (
    .a(al_b671fee2[4]),
    .b(al_45d9e18e[4]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_c325b022[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*C))+B*A*~((D*C))+~(B)*A*(D*C)+B*A*(D*C))"),
    .INIT(16'haccc))
    al_59a5b1c8 (
    .a(al_b671fee2[4]),
    .b(al_9892447e[4]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_1a25e1aa[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((D*~C))+B*A*~((D*~C))+~(B)*A*(D*~C)+B*A*(D*~C))"),
    .INIT(16'hcacc))
    al_50133ee1 (
    .a(al_b671fee2[4]),
    .b(al_c5e4c82d[4]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_6f7a76fc[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A)*~((~D*~C))+B*A*~((~D*~C))+~(B)*A*(~D*~C)+B*A*(~D*~C))"),
    .INIT(16'hccca))
    al_13bd720f (
    .a(al_b671fee2[4]),
    .b(al_89ad3a7d[4]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_2497ff95[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0aaaaff00))
    al_7220e142 (
    .a(al_c325b022[4]),
    .b(al_1a25e1aa[4]),
    .c(al_6f7a76fc[4]),
    .d(al_2497ff95[4]),
    .e(al_b1a73cf[0]),
    .f(al_b1a73cf[1]),
    .o(al_5b784e0e[4]));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    al_dfd625a4 (
    .a(al_a6bfe69c),
    .b(al_a09b37ae),
    .c(al_ef35f7b6[32]),
    .d(al_ef35f7b6[33]),
    .o(al_d271b0a3));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    al_5a12f7d1 (
    .a(al_263ba241),
    .b(al_50bc0ffd),
    .c(al_ef35f7b6[36]),
    .d(al_ef35f7b6[37]),
    .o(al_b537e59c));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*(D@C))"),
    .INIT(16'h0220))
    al_709f7cfe (
    .a(al_b537e59c),
    .b(al_4ee2ea2f),
    .c(al_440bddc2),
    .d(al_ef35f7b6[24]),
    .o(al_6df2ab59));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_74274fae (
    .a(al_65e4d4e0),
    .b(al_321810b0),
    .c(al_82001be8),
    .d(al_9941ff24[1]),
    .e(al_9941ff24[0]),
    .o(al_759a1829));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9a5528ab (
    .a(init_calib_complete),
    .b(al_6896ad14),
    .o(al_f7a41bbb));
  AL_MAP_LUT4 #(
    .EQN("(A*(~(B)*~(C)*~(D)+B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D+~(B)*C*D))"),
    .INIT(16'h282a))
    al_45447982 (
    .a(al_edebd92e),
    .b(al_9d2be50d[0]),
    .c(al_9d2be50d[1]),
    .d(al_530cb84f),
    .o(al_a57e41b7));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_f3df2499 (
    .a(al_6896ad14),
    .b(al_12521532),
    .o(al_52d7a8c5));
  AL_MAP_LUT6 #(
    .EQN("(F*~(~E*~D*C*~B*A))"),
    .INIT(64'hffffffdf00000000))
    al_fb18f3b (
    .a(al_65e4d4e0),
    .b(al_321810b0),
    .c(al_82001be8),
    .d(al_9941ff24[1]),
    .e(al_9941ff24[0]),
    .f(al_52d7a8c5),
    .o(al_61f2ed17));
  AL_MAP_LUT6 #(
    .EQN("(~((C*B*A))*D*~(E)*~(F)+~((C*B*A))*~(D)*E*~(F)+(C*B*A)*~(D)*E*~(F)+~((C*B*A))*D*E*~(F)+(C*B*A)*D*E*~(F)+~((C*B*A))*D*~(E)*F+~((C*B*A))*~(D)*E*F+~((C*B*A))*D*E*F)"),
    .INIT(64'h7f7f7f00ffff7f00))
    al_714c7ab9 (
    .a(al_a639b152),
    .b(al_386e051a),
    .c(al_6df2ab59),
    .d(al_759a1829),
    .e(al_61f2ed17),
    .f(al_1549e910),
    .o(al_f7d43aab));
  AL_MAP_LUT5 #(
    .EQN("(~D*C*~(E*~(B*A)))"),
    .INIT(32'h008000f0))
    al_b22e1865 (
    .a(al_58fb4752[3]),
    .b(al_58fb4752[4]),
    .c(al_f7a41bbb),
    .d(al_9d2be50d[0]),
    .e(al_12521532),
    .o(al_a7d66e26));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*B*~(E*A)))"),
    .INIT(32'h00bf003f))
    al_556e6a7f (
    .a(al_c088e9dc),
    .b(al_9d2be50d[0]),
    .c(al_9d2be50d[1]),
    .d(al_9d2be50d[2]),
    .e(al_c360bf4c[3]),
    .o(al_fc5dd8f9));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    al_801f8246 (
    .a(al_afc586c3),
    .b(al_6e8781e4),
    .c(al_ef35f7b6[29]),
    .o(al_a59a1785));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(D*~(~F*~(~C*~(E*~A)))))"),
    .INIT(64'h0033003331333033))
    al_e7ee04e3 (
    .a(al_f7d43aab),
    .b(al_a57e41b7),
    .c(al_a7d66e26),
    .d(al_fc5dd8f9),
    .e(al_9d2be50d[0]),
    .f(al_9d2be50d[1]),
    .o(al_7db277fb[0]));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*(E@D))"),
    .INIT(32'h00808000))
    al_23c7293 (
    .a(al_a59a1785),
    .b(al_d271b0a3),
    .c(al_6d82e9d5),
    .d(al_dc12b1d7),
    .e(al_ef35f7b6[25]),
    .o(al_a639b152));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    al_f27c93a1 (
    .a(al_4c7c6ba3),
    .b(al_d1e349fb),
    .c(al_ef35f7b6[26]),
    .d(al_ef35f7b6[27]),
    .o(al_f9cc5188));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*(D@C))"),
    .INIT(16'h0220))
    al_40033c4c (
    .a(al_f9cc5188),
    .b(al_5ea47e0d),
    .c(al_5fff4931),
    .d(al_ef35f7b6[28]),
    .o(al_386e051a));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*~(C*B*A))"),
    .INIT(64'h000000007f000000))
    al_644e80bb (
    .a(al_a639b152),
    .b(al_386e051a),
    .c(al_6df2ab59),
    .d(al_759a1829),
    .e(al_382cf878),
    .f(al_9d2be50d[2]),
    .o(al_7a15bb7a));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*~A))*~(B)+D*(C*~A)*~(B)+~(D)*(C*~A)*B+D*(C*~A)*B)"),
    .INIT(16'h8cbf))
    al_82eb2a8b (
    .a(al_c088e9dc),
    .b(al_9d2be50d[0]),
    .c(al_c360bf4c[3]),
    .d(al_4c58e022),
    .o(al_cc5fd2c8));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfc0faa00fc00aa00))
    al_86d27631 (
    .a(al_cc5fd2c8),
    .b(al_c088e9dc),
    .c(al_9d2be50d[0]),
    .d(al_9d2be50d[1]),
    .e(al_9d2be50d[2]),
    .f(al_530cb84f),
    .o(al_d244c645));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~A*~(~E*D*B))"),
    .INIT(32'hfafafefa))
    al_e2a55f4e (
    .a(al_7a15bb7a),
    .b(al_65bd6ac6),
    .c(al_d244c645),
    .d(al_382cf878),
    .e(al_9d2be50d[2]),
    .o(al_7db277fb[1]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    al_f5f0568f (
    .a(al_c088e9dc),
    .b(al_9d2be50d[0]),
    .c(al_c360bf4c[3]),
    .d(al_4c58e022),
    .o(al_e319e994));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfcf05500fcff5500))
    al_511e6261 (
    .a(al_e319e994),
    .b(al_c088e9dc),
    .c(al_9d2be50d[0]),
    .d(al_9d2be50d[1]),
    .e(al_9d2be50d[2]),
    .f(al_530cb84f),
    .o(al_7db277fb[2]));
  AL_MAP_LUT5 #(
    .EQN("((~B*A)*~(C)*~(D)*~(E)+(~B*A)*C*~(D)*~(E)+~((~B*A))*~(C)*D*~(E)+(~B*A)*~(C)*D*~(E)+~((~B*A))*C*~(D)*E+(~B*A)*C*~(D)*E+~((~B*A))*~(C)*D*E+(~B*A)*~(C)*D*E+~((~B*A))*C*D*E+(~B*A)*C*D*E)"),
    .INIT(32'hfff00f22))
    al_37dbf1eb (
    .a(al_8e6a6170),
    .b(al_fc44176c),
    .c(al_d51c2ed1),
    .d(al_10aff3dd[0]),
    .e(al_10aff3dd[1]),
    .o(al_4795b95a[0]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(~C*B*A))"),
    .INIT(16'hff08))
    al_113e5cc2 (
    .a(al_8e6a6170),
    .b(al_fc44176c),
    .c(al_10aff3dd[0]),
    .d(al_10aff3dd[1]),
    .o(al_4795b95a[1]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_5b568e25 (
    .a(al_c906bdb),
    .b(al_5a31c994),
    .c(al_56998d64),
    .o(al_3f4770be));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_b990f294 (
    .a(al_424bd4b9),
    .b(al_5a31c994),
    .c(al_56998d64),
    .o(al_509bee50));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_b96cfcaf (
    .a(al_802e0d75),
    .b(al_5a31c994),
    .c(al_56998d64),
    .o(al_3ec9b0d6));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_4c507cd8 (
    .a(al_cf11b78b[3]),
    .b(al_9d2be50d[0]),
    .c(al_9d2be50d[1]),
    .d(al_9d2be50d[2]),
    .e(al_898823b1),
    .o(al_5a31c994));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_85f8f86e (
    .a(al_2010f91b),
    .b(al_5a31c994),
    .c(al_56998d64),
    .o(al_eedba0b4));
  AL_DFF_0 al_ae98fa18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2af0d594),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_dd965664));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    al_3a0f78a9 (
    .a(al_7a15bb7a),
    .b(al_dd965664),
    .c(al_4c58e022),
    .o(al_2af0d594));
  AL_DFF_0 al_ce3c31e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f6114766[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_1a411806));
  AL_DFF_0 al_b0501b03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f6114766[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_6ea52063));
  AL_DFF_0 al_c5afcd1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f6114766[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_4d29fbf3));
  AL_DFF_0 al_a2d79ae0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f6114766[3]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_f2c5bff2));
  AL_DFF_0 al_71ecae42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f6114766[4]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_862761d2));
  AL_DFF_0 al_af396c2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a8314aee[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fb5f7a37));
  AL_DFF_0 al_9a76bc0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a8314aee[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_cc48041b));
  AL_DFF_0 al_6d936a16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a8314aee[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_cd905f33));
  AL_DFF_0 al_c192029e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a8314aee[3]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3151fa0));
  AL_DFF_0 al_b319aaf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff167b71[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_a879fe30));
  AL_DFF_0 al_a7cea116 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff167b71[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_bed6ed0d));
  AL_DFF_0 al_f80a14c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff167b71[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_8fadd979));
  AL_DFF_0 al_ee9306fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff167b71[3]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_28335c6e));
  AL_DFF_0 al_43796a92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_74d1b04e[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_5134abf1));
  AL_DFF_0 al_40845320 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_74d1b04e[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_d7e366bb));
  AL_DFF_0 al_8c26c73e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_74d1b04e[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_e8c2a90e));
  AL_DFF_0 al_1b3a698d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_74d1b04e[3]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_dd1e54e7));
  AL_DFF_0 al_e1da9286 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9d7bf9ff[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_824b4372));
  AL_DFF_0 al_8a140d92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9d7bf9ff[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_748a22bd));
  AL_DFF_0 al_1efbe077 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9d7bf9ff[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_6bd11777));
  AL_DFF_0 al_b2aa23de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9d7bf9ff[3]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_19255c36));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_5fe435f9 (
    .a(al_9d2be50d[0]),
    .b(al_9d2be50d[1]),
    .c(al_9d2be50d[2]),
    .o(al_a26ecd1c));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_6f88d3f6 (
    .a(al_a26ecd1c),
    .b(al_ef35f7b6[0]),
    .c(al_ef35f7b6[1]),
    .o(al_424bd4b9));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_485d849 (
    .a(al_424bd4b9),
    .b(al_c360bf4c[3]),
    .o(al_cce019));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_10695743 (
    .a(al_cce019),
    .b(al_a879fe30),
    .c(al_bed6ed0d),
    .d(al_8fadd979),
    .e(al_28335c6e),
    .f(al_6f5534a0),
    .o(al_ff167b71[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_d0df3865 (
    .a(al_cce019),
    .b(al_a879fe30),
    .c(al_6f5534a0),
    .o(al_ff167b71[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_64dd3ece (
    .a(al_cce019),
    .b(al_a879fe30),
    .c(al_bed6ed0d),
    .d(al_6f5534a0),
    .o(al_ff167b71[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_e294d786 (
    .a(al_cce019),
    .b(al_a879fe30),
    .c(al_bed6ed0d),
    .d(al_8fadd979),
    .e(al_6f5534a0),
    .o(al_ff167b71[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_76ec3733 (
    .a(al_a26ecd1c),
    .b(al_ef35f7b6[0]),
    .c(al_ef35f7b6[1]),
    .o(al_802e0d75));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_123cd809 (
    .a(al_802e0d75),
    .b(al_c360bf4c[3]),
    .o(al_31bcb2f7));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_229eff30 (
    .a(al_31bcb2f7),
    .b(al_5134abf1),
    .c(al_d7e366bb),
    .d(al_e8c2a90e),
    .e(al_dd1e54e7),
    .f(al_f1c7f7af),
    .o(al_74d1b04e[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_a208a457 (
    .a(al_31bcb2f7),
    .b(al_5134abf1),
    .c(al_f1c7f7af),
    .o(al_74d1b04e[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_d841d122 (
    .a(al_31bcb2f7),
    .b(al_5134abf1),
    .c(al_d7e366bb),
    .d(al_f1c7f7af),
    .o(al_74d1b04e[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_23639d04 (
    .a(al_31bcb2f7),
    .b(al_5134abf1),
    .c(al_d7e366bb),
    .d(al_e8c2a90e),
    .e(al_f1c7f7af),
    .o(al_74d1b04e[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_3aa91860 (
    .a(al_a26ecd1c),
    .b(al_ef35f7b6[0]),
    .c(al_ef35f7b6[1]),
    .o(al_2010f91b));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_786fd53d (
    .a(al_2010f91b),
    .b(al_c360bf4c[3]),
    .o(al_b887382e));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_f9a2df13 (
    .a(al_b887382e),
    .b(al_824b4372),
    .c(al_748a22bd),
    .d(al_6bd11777),
    .e(al_19255c36),
    .f(al_cf38d855),
    .o(al_9d7bf9ff[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_1c46400 (
    .a(al_b887382e),
    .b(al_824b4372),
    .c(al_cf38d855),
    .o(al_9d7bf9ff[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_d2b3a674 (
    .a(al_b887382e),
    .b(al_824b4372),
    .c(al_748a22bd),
    .d(al_cf38d855),
    .o(al_9d7bf9ff[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_50bf5fdb (
    .a(al_b887382e),
    .b(al_824b4372),
    .c(al_748a22bd),
    .d(al_6bd11777),
    .e(al_cf38d855),
    .o(al_9d7bf9ff[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_45cbde2c (
    .a(al_a26ecd1c),
    .b(al_ef35f7b6[0]),
    .c(al_ef35f7b6[1]),
    .o(al_c906bdb));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9f334e8a (
    .a(al_c906bdb),
    .b(al_c360bf4c[3]),
    .o(al_da7de1b7));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E@(~F*~D*~C*~B)))"),
    .INIT(64'h5555000055540001))
    al_e91f5861 (
    .a(al_da7de1b7),
    .b(al_fb5f7a37),
    .c(al_cc48041b),
    .d(al_cd905f33),
    .e(al_3151fa0),
    .f(al_63204f4),
    .o(al_a8314aee[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    al_8544ac44 (
    .a(al_da7de1b7),
    .b(al_fb5f7a37),
    .c(al_63204f4),
    .o(al_a8314aee[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(~D*~B)))"),
    .INIT(16'h5041))
    al_f3fdc351 (
    .a(al_da7de1b7),
    .b(al_fb5f7a37),
    .c(al_cc48041b),
    .d(al_63204f4),
    .o(al_a8314aee[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(D@(~E*~C*~B)))"),
    .INIT(32'h55005401))
    al_28fd42f (
    .a(al_da7de1b7),
    .b(al_fb5f7a37),
    .c(al_cc48041b),
    .d(al_cd905f33),
    .e(al_63204f4),
    .o(al_a8314aee[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_2e3ac9d2 (
    .a(al_ff167b71[3]),
    .b(al_ff167b71[0]),
    .c(al_ff167b71[1]),
    .d(al_ff167b71[2]),
    .o(al_251b6a5[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_d2290915 (
    .a(al_74d1b04e[3]),
    .b(al_74d1b04e[0]),
    .c(al_74d1b04e[1]),
    .d(al_74d1b04e[2]),
    .o(al_251b6a5[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_adc9c3a6 (
    .a(al_9d7bf9ff[3]),
    .b(al_9d7bf9ff[0]),
    .c(al_9d7bf9ff[1]),
    .d(al_9d7bf9ff[2]),
    .o(al_251b6a5[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_2d660cdd (
    .a(al_a8314aee[3]),
    .b(al_a8314aee[0]),
    .c(al_a8314aee[1]),
    .d(al_a8314aee[2]),
    .o(al_251b6a5[0]));
  AL_DFF_0 al_3cc3c2d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_251b6a5[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_63204f4));
  AL_DFF_0 al_fed05e12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_251b6a5[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f5534a0));
  AL_DFF_0 al_23c2ba7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_251b6a5[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1c7f7af));
  AL_DFF_0 al_be58b012 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_251b6a5[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf38d855));
  AL_DFF_0 al_ad2da7c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ffc3eff4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c1c29ee));
  AL_DFF_0 al_322b0c9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[24]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2f7a19ec));
  AL_DFF_0 al_5e0d281b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[25]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_41c51f8));
  AL_DFF_0 al_5329199c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[26]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b169d8ec));
  AL_DFF_0 al_fe0edfb6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[27]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c4782d2));
  AL_DFF_0 al_6e45321b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[28]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3d92dfa6));
  AL_DFF_0 al_7db12f17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[29]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_49679814));
  AL_DFF_0 al_49cb3e12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[30]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_884f3fa8));
  AL_DFF_0 al_c6def0ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[31]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_13d7dde4));
  AL_DFF_0 al_576121f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[32]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b63d0e11));
  AL_DFF_0 al_11aa4253 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[33]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2819b010));
  AL_DFF_0 al_1f94ace9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[34]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_c64ad91c));
  AL_DFF_0 al_3d727427 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[35]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_c81413d1));
  AL_DFF_0 al_22221731 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[36]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_4aecdf04));
  AL_DFF_0 al_f1ff6d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[37]),
    .en(al_3f4770be),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2024cd4b));
  AL_DFF_0 al_8dbadb4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_526ace65),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d99a742));
  AL_DFF_0 al_ca1071e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[24]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_d301de48));
  AL_DFF_0 al_1db7f656 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[25]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_ce2e94ee));
  AL_DFF_0 al_e7232016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[26]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_44e6dfe9));
  AL_DFF_0 al_fff3d7c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[27]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b091346b));
  AL_DFF_0 al_54940863 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[28]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_e4f5dc3f));
  AL_DFF_0 al_fe521d0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[29]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_c2e0ff4));
  AL_DFF_0 al_3b8ebe3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[30]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_91bd4a18));
  AL_DFF_0 al_a5eadb34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[31]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_4c19e182));
  AL_DFF_0 al_21e2c40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[32]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_46d55200));
  AL_DFF_0 al_cf11a9cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[33]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_98c513dd));
  AL_DFF_0 al_8e0c86e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[34]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_5ae0756d));
  AL_DFF_0 al_5ff83d4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[35]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_5f6a6401));
  AL_DFF_0 al_28736b7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[36]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_dcf6b718));
  AL_DFF_0 al_a9e1f46c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[37]),
    .en(al_509bee50),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_4e84d779));
  AL_DFF_0 al_e50c95fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3514085d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1001936c));
  AL_DFF_0 al_4d4e54ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[24]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_963a39c1));
  AL_DFF_0 al_197c32bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[25]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_bc5117fe));
  AL_DFF_0 al_2432ae52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[26]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_92d8fd60));
  AL_DFF_0 al_d7dacb1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[27]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_126719a0));
  AL_DFF_0 al_550f41b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[28]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_e8289617));
  AL_DFF_0 al_80c4a66d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[29]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_bc7b13ca));
  AL_DFF_0 al_140f9bb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[30]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_1b5b7fb8));
  AL_DFF_0 al_1c9495b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[31]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_316deb29));
  AL_DFF_0 al_ba30a8b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[32]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7e44c8d5));
  AL_DFF_0 al_3150fe37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[33]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_74066232));
  AL_DFF_0 al_fc2eeab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[34]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7eff70ba));
  AL_DFF_0 al_f2dd49c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[35]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9bbade9e));
  AL_DFF_0 al_9b1f88c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[36]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_91941257));
  AL_DFF_0 al_80941e84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[37]),
    .en(al_3ec9b0d6),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_df5d8efd));
  AL_DFF_0 al_ead02cfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_270372c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c61f1e9a));
  AL_DFF_0 al_79e9031d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[24]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3f2ddb8a));
  AL_DFF_0 al_ca68c870 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[25]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_8fd7f3b8));
  AL_DFF_0 al_6ec18378 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[26]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7059c89d));
  AL_DFF_0 al_2474eb57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[27]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_ed48bce4));
  AL_DFF_0 al_622527d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[28]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_6b5d2018));
  AL_DFF_0 al_45462fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[29]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7564e3b0));
  AL_DFF_0 al_6ae70728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[30]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3f998e21));
  AL_DFF_0 al_2ebbd834 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[31]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2115cf8f));
  AL_DFF_0 al_cadb4c8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[32]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_f7549f58));
  AL_DFF_0 al_30ddc37e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[33]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_f3529ba5));
  AL_DFF_0 al_29691bd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[34]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_a0f5de0d));
  AL_DFF_0 al_d1ba9df7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[35]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3bcdd651));
  AL_DFF_0 al_94e54eed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[36]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_47aa4bf9));
  AL_DFF_0 al_fc682ebb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[37]),
    .en(al_eedba0b4),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_5758806f));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_222d70e3 (
    .a(al_424bd4b9),
    .b(al_5a31c994),
    .c(al_9d99a742),
    .d(al_56998d64),
    .e(al_4dd68878),
    .o(al_526ace65));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_e15299ff (
    .a(al_c906bdb),
    .b(al_5a31c994),
    .c(al_5c1c29ee),
    .d(al_56998d64),
    .e(al_4dd68878),
    .o(al_ffc3eff4));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_d15aa9bb (
    .a(al_2010f91b),
    .b(al_5a31c994),
    .c(al_c61f1e9a),
    .d(al_56998d64),
    .e(al_4dd68878),
    .o(al_270372c));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~A*~(C*~B)))"),
    .INIT(32'h000000ba))
    al_b3d83db3 (
    .a(al_802e0d75),
    .b(al_5a31c994),
    .c(al_1001936c),
    .d(al_56998d64),
    .e(al_4dd68878),
    .o(al_3514085d));
  AL_DFF_0 al_7f56392a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71faa803[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56998d64));
  AL_DFF_0 al_ebfd710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c4fa309[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_c28589ac));
  AL_DFF_0 al_1a6af1d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9a0a15b5),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_198de9a1));
  AL_MAP_LUT6 #(
    .EQN("(~C*~(~D*~(~F*~E*B*A)))"),
    .INIT(64'h0f000f000f000f08))
    al_c41cc021 (
    .a(al_8e6a6170),
    .b(al_238af9ad),
    .c(al_d51c2ed1),
    .d(al_198de9a1),
    .e(al_10aff3dd[0]),
    .f(al_10aff3dd[1]),
    .o(al_9a0a15b5));
  AL_DFF_0 al_5fbd11c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_68e89a39),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cf11b78b[3]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_ad9843a (
    .a(al_6896ad14),
    .b(al_d149d704),
    .c(al_9d2be50d[0]),
    .d(al_9d2be50d[1]),
    .e(al_9d2be50d[2]),
    .o(al_68e89a39));
  AL_DFF_0 al_3421cfdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_93070309),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbeafa67[6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    al_daa329fc (
    .a(al_7a15bb7a),
    .b(al_cbeafa67[6]),
    .c(al_ef35f7b6[2]),
    .d(al_4dd68878),
    .o(al_93070309));
  AL_DFF_0 al_e4657a06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_4ed70d21[0]));
  AL_DFF_0 al_db46b6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_4ed70d21[1]));
  AL_DFF_0 al_f50aef7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_d76fa964[6]));
  AL_DFF_0 al_8565099a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7db277fb[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9d2be50d[0]));
  AL_DFF_0 al_8e0db69a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7db277fb[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9d2be50d[1]));
  AL_DFF_0 al_cc5a9539 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7db277fb[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9d2be50d[2]));
  AL_DFF_0 al_43ad039 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4795b95a[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_10aff3dd[0]));
  AL_DFF_0 al_60d61bb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4795b95a[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_10aff3dd[1]));
  AL_DFF_0 al_fbbeaf5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2497ff95[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89ad3a7d[0]));
  AL_DFF_0 al_268952db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2497ff95[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89ad3a7d[1]));
  AL_DFF_0 al_1033f88d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2497ff95[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89ad3a7d[2]));
  AL_DFF_0 al_9fa620a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2497ff95[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89ad3a7d[3]));
  AL_DFF_0 al_eca57e04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2497ff95[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89ad3a7d[4]));
  AL_DFF_0 al_22375e7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c325b022[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45d9e18e[0]));
  AL_DFF_0 al_d6479572 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c325b022[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45d9e18e[1]));
  AL_DFF_0 al_b658168d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c325b022[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45d9e18e[2]));
  AL_DFF_0 al_745e738f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c325b022[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45d9e18e[3]));
  AL_DFF_0 al_4e94cbb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c325b022[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45d9e18e[4]));
  AL_DFF_0 al_bea51882 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6f7a76fc[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5e4c82d[0]));
  AL_DFF_0 al_5ed6265e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6f7a76fc[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5e4c82d[1]));
  AL_DFF_0 al_f48f1a88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6f7a76fc[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5e4c82d[2]));
  AL_DFF_0 al_4c35ca8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6f7a76fc[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5e4c82d[3]));
  AL_DFF_0 al_91078e8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6f7a76fc[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5e4c82d[4]));
  AL_DFF_0 al_84e81e37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a25e1aa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9892447e[0]));
  AL_DFF_0 al_7b3e601e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a25e1aa[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9892447e[1]));
  AL_DFF_0 al_633d4ca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a25e1aa[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9892447e[2]));
  AL_DFF_0 al_830e9af5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a25e1aa[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9892447e[3]));
  AL_DFF_0 al_228479db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a25e1aa[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9892447e[4]));
  AL_DFF_0 al_2ba55e6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba0505cb[3]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7054a209[3]));
  AL_DFF_0 al_fdd7f5e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba0505cb[4]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7054a209[4]));
  AL_DFF_0 al_f5b086f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba0505cb[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7054a209[0]));
  AL_DFF_0 al_90907e9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba0505cb[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7054a209[1]));
  AL_DFF_0 al_83cb301e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba0505cb[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_7054a209[2]));
  AL_DFF_0 al_6556bc7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[0]));
  AL_DFF_0 al_ddbfee29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[1]));
  AL_DFF_0 al_d02927b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[2]));
  AL_DFF_0 al_21d39dc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[11]));
  AL_DFF_0 al_55421e18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[12]));
  AL_DFF_0 al_1b5a1f77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[13]));
  AL_DFF_0 al_3092364e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[14]));
  AL_DFF_0 al_9973a77c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[15]));
  AL_DFF_0 al_f0a27c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[16]));
  AL_DFF_0 al_4740c96d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[17]));
  AL_DFF_0 al_d44c1ffd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[24]));
  AL_DFF_0 al_14476f1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[25]));
  AL_DFF_0 al_d6b7a2e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[26]));
  AL_DFF_0 al_fca9e724 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[27]));
  AL_DFF_0 al_98e49513 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[28]));
  AL_DFF_0 al_d2f5df57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[29]));
  AL_DFF_0 al_cfc5b4ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[30]));
  AL_DFF_0 al_8f1d5574 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[31]));
  AL_DFF_0 al_44124080 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[32]));
  AL_DFF_0 al_d1d442df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[33]));
  AL_DFF_0 al_616d72eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[34]));
  AL_DFF_0 al_faab6e47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[35]));
  AL_DFF_0 al_a19f98b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[36]));
  AL_DFF_0 al_77f36fa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[37]));
  AL_DFF_0 al_19dd3733 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[44]));
  AL_DFF_0 al_5c60ce6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[45]));
  AL_DFF_0 al_de8fbf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_786f2a14[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef35f7b6[46]));
  AL_DFF_0 al_7132dce1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[0]));
  AL_DFF_0 al_aa7e20f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[1]));
  AL_DFF_0 al_77747a73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[2]));
  AL_DFF_0 al_5ca53269 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[11]));
  AL_DFF_0 al_41ecf4f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[12]));
  AL_DFF_0 al_7bd91581 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[13]));
  AL_DFF_0 al_a989bd2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[14]));
  AL_DFF_0 al_d3f024a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[15]));
  AL_DFF_0 al_e60fa356 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[16]));
  AL_DFF_0 al_384f454c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[17]));
  AL_DFF_0 al_ea069cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[24]));
  AL_DFF_0 al_6555d9c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[25]));
  AL_DFF_0 al_e1e36854 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[26]));
  AL_DFF_0 al_61f5a813 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[27]));
  AL_DFF_0 al_bbb765cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[28]));
  AL_DFF_0 al_e21d1730 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[29]));
  AL_DFF_0 al_835f5f0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[30]));
  AL_DFF_0 al_2511d03a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[31]));
  AL_DFF_0 al_ec7fb03d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[32]));
  AL_DFF_0 al_453184cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[33]));
  AL_DFF_0 al_15e1b6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[34]));
  AL_DFF_0 al_ae4786b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[35]));
  AL_DFF_0 al_b1f01e5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[36]));
  AL_DFF_0 al_c554de8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[37]));
  AL_DFF_0 al_ccd7e764 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[44]));
  AL_DFF_0 al_39e626fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[45]));
  AL_DFF_0 al_15789529 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_f001c0eb[0]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_3c07b31a[46]));
  AL_DFF_0 al_8cc5ac49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[0]));
  AL_DFF_0 al_9e951d40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[1]));
  AL_DFF_0 al_d47e1e2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[2]));
  AL_DFF_0 al_ffdb003 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[11]));
  AL_DFF_0 al_f40b5875 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[12]));
  AL_DFF_0 al_e1d6378b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[13]));
  AL_DFF_0 al_7bd1d88e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[14]));
  AL_DFF_0 al_9ff2f8d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[15]));
  AL_DFF_0 al_6c383fcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[16]));
  AL_DFF_0 al_c44eb6da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[17]));
  AL_DFF_0 al_a124ae8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[24]));
  AL_DFF_0 al_63d5597f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[25]));
  AL_DFF_0 al_928cacc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[26]));
  AL_DFF_0 al_6c22bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[27]));
  AL_DFF_0 al_e77c7797 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[28]));
  AL_DFF_0 al_a83e668d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[29]));
  AL_DFF_0 al_9cceb6e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[30]));
  AL_DFF_0 al_8f06360d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[31]));
  AL_DFF_0 al_50b381ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[32]));
  AL_DFF_0 al_f098fda1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[33]));
  AL_DFF_0 al_d8ccd401 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[34]));
  AL_DFF_0 al_3d0423ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[35]));
  AL_DFF_0 al_cff06948 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[36]));
  AL_DFF_0 al_af6a79e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[37]));
  AL_DFF_0 al_81d5a612 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[44]));
  AL_DFF_0 al_202bdaf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[45]));
  AL_DFF_0 al_7124d97f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_f001c0eb[1]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_fbcce8b0[46]));
  AL_DFF_0 al_fa9ec201 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[0]));
  AL_DFF_0 al_348ccb5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[1]));
  AL_DFF_0 al_eadc4bf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[2]));
  AL_DFF_0 al_23e38e90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[11]));
  AL_DFF_0 al_ce19996f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[12]));
  AL_DFF_0 al_5803d5e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[13]));
  AL_DFF_0 al_a2bb4d9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[14]));
  AL_DFF_0 al_2088e866 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[15]));
  AL_DFF_0 al_9d3a8fd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[16]));
  AL_DFF_0 al_5130b66e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[17]));
  AL_DFF_0 al_92417236 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[24]));
  AL_DFF_0 al_35d87eae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[25]));
  AL_DFF_0 al_a1ee9419 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[26]));
  AL_DFF_0 al_3cf819de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[27]));
  AL_DFF_0 al_600b6ac1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[28]));
  AL_DFF_0 al_5cb657d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[29]));
  AL_DFF_0 al_7cdec05a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[30]));
  AL_DFF_0 al_effdafb6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[31]));
  AL_DFF_0 al_23bff2b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[32]));
  AL_DFF_0 al_89033031 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[33]));
  AL_DFF_0 al_eb662a12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[34]));
  AL_DFF_0 al_cd5497ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[35]));
  AL_DFF_0 al_9ccb8e78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[36]));
  AL_DFF_0 al_926b7901 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[37]));
  AL_DFF_0 al_52cd224 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[44]));
  AL_DFF_0 al_a27b8010 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[45]));
  AL_DFF_0 al_d263fcc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_f001c0eb[2]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2422b44d[46]));
  AL_DFF_0 al_87786687 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[5]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[0]));
  AL_DFF_0 al_9df3f1dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[3]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[1]));
  AL_DFF_0 al_c08c745a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[4]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[2]));
  AL_DFF_0 al_4a086558 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[6]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[11]));
  AL_DFF_0 al_9f51d970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[7]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[12]));
  AL_DFF_0 al_80082e4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[8]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[13]));
  AL_DFF_0 al_699fabdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[9]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[14]));
  AL_DFF_0 al_1ff04b09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[10]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[15]));
  AL_DFF_0 al_21d21c55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[11]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[16]));
  AL_DFF_0 al_18b3ff1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[12]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[17]));
  AL_DFF_0 al_64bc2af8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[13]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[24]));
  AL_DFF_0 al_356fa8bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[14]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[25]));
  AL_DFF_0 al_d443226d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[15]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[26]));
  AL_DFF_0 al_592e532d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[16]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[27]));
  AL_DFF_0 al_888610f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[17]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[28]));
  AL_DFF_0 al_9aa2db47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[18]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[29]));
  AL_DFF_0 al_423d0573 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[19]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[30]));
  AL_DFF_0 al_7bbe926c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[20]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[31]));
  AL_DFF_0 al_fc91a138 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[21]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[32]));
  AL_DFF_0 al_72000ca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[22]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[33]));
  AL_DFF_0 al_204951ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[23]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[34]));
  AL_DFF_0 al_a45c67b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[24]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[35]));
  AL_DFF_0 al_dc235ec1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[25]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[36]));
  AL_DFF_0 al_c962bd3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_58fb4752[26]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[37]));
  AL_DFF_0 al_b4978c59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[44]));
  AL_DFF_0 al_f1588e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[45]));
  AL_DFF_0 al_3a2f643a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(al_f001c0eb[3]),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_9c80d3c6[46]));
  AL_DFF_0 al_a2427aa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e11b20ed[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b1a73cf[0]));
  AL_DFF_0 al_f3d8b60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e11b20ed[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b1a73cf[1]));
  AL_DFF_0 al_1cf46c5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1373d93[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_1124d2df[0]));
  AL_DFF_0 al_159417d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a1373d93[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_1124d2df[1]));
  AL_DFF_0 al_e5d91fca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[0]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd768853[0]));
  AL_DFF_0 al_2f2eeecf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[1]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd768853[1]));
  AL_DFF_0 al_ce25a088 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[2]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd768853[2]));
  AL_DFF_0 al_ea001341 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[3]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd768853[3]));
  AL_DFF_0 al_24b67d4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[4]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd768853[4]));
  AL_DFF_0 al_7165900f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[0]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec54698[0]));
  AL_DFF_0 al_5cb5ec3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[1]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec54698[1]));
  AL_DFF_0 al_11d7303b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[2]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec54698[2]));
  AL_DFF_0 al_fd3c3aa3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[3]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec54698[3]));
  AL_DFF_0 al_166ef66b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[4]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec54698[4]));
  AL_DFF_0 al_a63ebb50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[0]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ffdc699f[0]));
  AL_DFF_0 al_10694171 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[1]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ffdc699f[1]));
  AL_DFF_0 al_3dd42822 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[2]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ffdc699f[2]));
  AL_DFF_0 al_81b48b70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[3]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ffdc699f[3]));
  AL_DFF_0 al_26d55608 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[4]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ffdc699f[4]));
  AL_DFF_0 al_e3aab822 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[0]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1974c03[0]));
  AL_DFF_0 al_bdfd3741 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[1]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1974c03[1]));
  AL_DFF_0 al_33439642 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[2]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1974c03[2]));
  AL_DFF_0 al_ad19d53a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[3]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1974c03[3]));
  AL_DFF_0 al_83f80465 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b784e0e[4]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1974c03[4]));
  AL_DFF_0 al_8553d7df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_68f1a7a7[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_a196b5f4[0]));
  AL_DFF_0 al_168d40b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_68f1a7a7[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_a196b5f4[1]));
  AL_DFF_0 al_e9597224 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_696c7934[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b25d0e99[0]));
  AL_DFF_0 al_b078dcee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_696c7934[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b25d0e99[1]));
  AL_DFF_0 al_e4fa35b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_696c7934[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b25d0e99[2]));
  AL_DFF_0 al_6b8785f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_696c7934[3]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_b25d0e99[3]));
  AL_DFF_0 al_28a98264 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[0]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[0]));
  AL_DFF_0 al_a9e9ddd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[1]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[1]));
  AL_DFF_0 al_b92c6e36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[2]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[2]));
  AL_DFF_0 al_446bd96d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[11]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[11]));
  AL_DFF_0 al_48edc538 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[12]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[12]));
  AL_DFF_0 al_85fe7b60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[13]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[13]));
  AL_DFF_0 al_2df3ec22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[14]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[14]));
  AL_DFF_0 al_4cc7f662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[15]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[15]));
  AL_DFF_0 al_2fc897b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[16]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[16]));
  AL_DFF_0 al_e2614b36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[17]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[17]));
  AL_DFF_0 al_9c1bc2aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[44]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[44]));
  AL_DFF_0 al_cddbf882 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[45]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[45]));
  AL_DFF_0 al_fbfdc32a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[46]),
    .en(al_69c2ff54[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_974136cc[46]));
  AL_DFF_0 al_5dd7cfc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[0]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[0]));
  AL_DFF_0 al_8cee241a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[1]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[1]));
  AL_DFF_0 al_36387710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[2]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[2]));
  AL_DFF_0 al_74e2390c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[11]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[11]));
  AL_DFF_0 al_d220ffe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[12]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[12]));
  AL_DFF_0 al_3f1c5dc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[13]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[13]));
  AL_DFF_0 al_cf1e0e1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[14]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[14]));
  AL_DFF_0 al_1b011c99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[15]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[15]));
  AL_DFF_0 al_50b8938 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[16]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[16]));
  AL_DFF_0 al_4e953b2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[17]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[17]));
  AL_DFF_0 al_1007f926 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[44]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[44]));
  AL_DFF_0 al_5f20775c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[45]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[45]));
  AL_DFF_0 al_86b61a8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[46]),
    .en(al_69c2ff54[1]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea7bbd9[46]));
  AL_DFF_0 al_fbd7f7e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[0]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[0]));
  AL_DFF_0 al_3dbed882 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[1]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[1]));
  AL_DFF_0 al_42ea5b39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[2]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[2]));
  AL_DFF_0 al_99b5c261 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[11]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[11]));
  AL_DFF_0 al_bd21cb48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[12]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[12]));
  AL_DFF_0 al_abf01007 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[13]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[13]));
  AL_DFF_0 al_d2c743a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[14]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[14]));
  AL_DFF_0 al_70fb3bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[15]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[15]));
  AL_DFF_0 al_c42d372c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[16]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[16]));
  AL_DFF_0 al_ac4c3743 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[17]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[17]));
  AL_DFF_0 al_dde7ecdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[44]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[44]));
  AL_DFF_0 al_2593fdc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[45]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[45]));
  AL_DFF_0 al_e809e59b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[46]),
    .en(al_69c2ff54[2]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16b7523e[46]));
  AL_DFF_0 al_c6974391 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[0]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[0]));
  AL_DFF_0 al_93af710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[1]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[1]));
  AL_DFF_0 al_7e97241e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[2]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[2]));
  AL_DFF_0 al_78277917 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[11]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[11]));
  AL_DFF_0 al_4fafffb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[12]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[12]));
  AL_DFF_0 al_44645df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[13]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[13]));
  AL_DFF_0 al_41167f57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[14]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[14]));
  AL_DFF_0 al_940a83a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[15]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[15]));
  AL_DFF_0 al_f7e488a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[16]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[16]));
  AL_DFF_0 al_a13d8daf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[17]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[17]));
  AL_DFF_0 al_71afb3da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[44]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[44]));
  AL_DFF_0 al_cc0661c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[45]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[45]));
  AL_DFF_0 al_596de69a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef35f7b6[46]),
    .en(al_69c2ff54[3]),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f82ace94[46]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    al_1f3e294d (
    .a(al_7a15bb7a),
    .b(al_ef35f7b6[0]),
    .c(al_53bb123b[6]),
    .d(al_4dd68878),
    .o(al_965bd4e5));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    al_5e01c1d (
    .a(al_7a15bb7a),
    .b(al_ef35f7b6[1]),
    .c(al_53bb123b[7]),
    .d(al_4dd68878),
    .o(al_8954e1e7));
  AL_DFF_0 al_93488869 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_965bd4e5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53bb123b[6]));
  AL_DFF_0 al_94056225 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8954e1e7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53bb123b[7]));
  AL_DFF_0 al_632a6065 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f7dedc[3]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_553ae5af[3]));
  AL_DFF_0 al_2e8b31af (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f7dedc[4]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_553ae5af[4]));
  AL_DFF_0 al_32523093 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f7dedc[0]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_553ae5af[0]));
  AL_DFF_0 al_a701778c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f7dedc[1]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_553ae5af[1]));
  AL_DFF_0 al_3d68dac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f7dedc[2]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_553ae5af[2]));
  AL_DFF_0 al_fd665810 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[11]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2602b5cf[33]));
  AL_DFF_0 al_9a1a6245 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[12]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2602b5cf[34]));
  AL_DFF_0 al_3c25f60b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[13]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2602b5cf[35]));
  AL_DFF_0 al_15783271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[14]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2602b5cf[36]));
  AL_DFF_0 al_9dbf7298 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[15]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2602b5cf[37]));
  AL_DFF_0 al_ffd00f1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[16]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2602b5cf[38]));
  AL_DFF_0 al_63224183 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7040e81f[17]),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_2602b5cf[39]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8d47c0a (
    .i(al_a3c26eaf),
    .o(al_53334a6));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3736997 (
    .i(al_53334a6),
    .o(al_4dd68878));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*B*~(C)*D*E)"),
    .INIT(32'h0800fbcf))
    al_13612fe4 (
    .a(al_1a411806),
    .b(al_9d2be50d[0]),
    .c(al_9d2be50d[1]),
    .d(al_9d2be50d[2]),
    .e(al_7054a209[0]),
    .o(al_ba0505cb[0]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haacaa0aa))
    al_aa2124bb (
    .a(al_e6d81dbe[4]),
    .b(al_862761d2),
    .c(al_9d2be50d[0]),
    .d(al_9d2be50d[1]),
    .e(al_9d2be50d[2]),
    .o(al_ba0505cb[4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_625e4442 (
    .a(al_ba0505cb[4]),
    .b(al_ba0505cb[3]),
    .c(al_ba0505cb[2]),
    .d(al_ba0505cb[1]),
    .e(al_ba0505cb[0]),
    .o(al_e650be8a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~((F@E))+A*~(B)*~(C)*~(D)*~((F@E))+~(A)*B*~(C)*~(D)*~((F@E))+A*B*~(C)*~(D)*~((F@E))+~(A)*B*C*~(D)*~((F@E))+A*B*C*~(D)*~((F@E))+~(A)*~(B)*~(C)*D*~((F@E))+A*~(B)*~(C)*D*~((F@E))+A*B*~(C)*D*~((F@E))+~(A)*~(B)*C*D*~((F@E))+A*~(B)*C*D*~((F@E))+~(A)*B*C*D*~((F@E))+A*B*C*D*~((F@E))+A*B*~(C)*D*(F@E))"),
    .INIT(64'hfbcf08000800fbcf))
    al_eb2fa568 (
    .a(al_6ea52063),
    .b(al_9d2be50d[0]),
    .c(al_9d2be50d[1]),
    .d(al_9d2be50d[2]),
    .e(al_7054a209[0]),
    .f(al_7054a209[1]),
    .o(al_ba0505cb[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C@(~B*~A))"),
    .INIT(8'h1e))
    al_51bf6349 (
    .a(al_7054a209[0]),
    .b(al_7054a209[1]),
    .c(al_7054a209[2]),
    .o(al_d4f7298c));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55c55055))
    al_abf0a28d (
    .a(al_d4f7298c),
    .b(al_4d29fbf3),
    .c(al_9d2be50d[0]),
    .d(al_9d2be50d[1]),
    .e(al_9d2be50d[2]),
    .o(al_ba0505cb[2]));
  AL_MAP_LUT4 #(
    .EQN("~(D@(~C*~B*~A))"),
    .INIT(16'h01fe))
    al_d76efea3 (
    .a(al_7054a209[0]),
    .b(al_7054a209[1]),
    .c(al_7054a209[2]),
    .d(al_7054a209[3]),
    .o(al_b1a37b71));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55c55055))
    al_d7621819 (
    .a(al_b1a37b71),
    .b(al_f2c5bff2),
    .c(al_9d2be50d[0]),
    .d(al_9d2be50d[1]),
    .e(al_9d2be50d[2]),
    .o(al_ba0505cb[3]));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~C*~B*~A))"),
    .INIT(32'hfffe0001))
    al_e5ae444c (
    .a(al_7054a209[0]),
    .b(al_7054a209[1]),
    .c(al_7054a209[2]),
    .d(al_7054a209[3]),
    .e(al_7054a209[4]),
    .o(al_e6d81dbe[4]));
  AL_DFF_0 al_8e126ee9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e650be8a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_530cb84f));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_2fbf7423 (
    .a(al_3e56391),
    .b(al_1124d2df[0]),
    .o(al_a1373d93[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    al_88c1407b (
    .a(al_3e56391),
    .b(al_1124d2df[0]),
    .c(al_1124d2df[1]),
    .o(al_a1373d93[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_829aec37 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_a1373d93[0]),
    .d(al_a1373d93[1]),
    .o(al_ce2030ae));
  AL_DFF_0 al_dea7f7f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ce2030ae),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12521532));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5cd12496 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[5]),
    .c(al_5d3f410a[5]),
    .o(al_58fb4752[5]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_406b6d20 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[5]),
    .c(al_3c07b31a[0]),
    .o(al_388ebe26));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ceb609da (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[5]),
    .c(al_fbcce8b0[0]),
    .o(al_d6e945fd[0]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_afb924d4 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[5]),
    .c(al_2422b44d[0]),
    .o(al_48b96055));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_dd9ebfff (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[5]),
    .c(al_9c80d3c6[0]),
    .o(al_f152e67e[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_8c4986a (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_388ebe26),
    .d(al_48b96055),
    .e(al_d6e945fd[0]),
    .f(al_f152e67e[0]),
    .o(al_786f2a14[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3e4c14de (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[6]),
    .c(al_5d3f410a[6]),
    .o(al_58fb4752[6]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_5bd84e2f (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[6]),
    .c(al_3c07b31a[11]),
    .o(al_a96965a6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_20a0898f (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[6]),
    .c(al_fbcce8b0[11]),
    .o(al_d6e945fd[11]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_12d1cfc5 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[6]),
    .c(al_2422b44d[11]),
    .o(al_bb6dcd3));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b8917cb6 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[6]),
    .c(al_9c80d3c6[11]),
    .o(al_f152e67e[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_112f6cb0 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_a96965a6),
    .d(al_bb6dcd3),
    .e(al_d6e945fd[11]),
    .f(al_f152e67e[11]),
    .o(al_786f2a14[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_95fd014f (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[7]),
    .c(al_5d3f410a[7]),
    .o(al_58fb4752[7]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_699abddb (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[7]),
    .c(al_3c07b31a[12]),
    .o(al_d3f078c4));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d6815c9e (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[7]),
    .c(al_fbcce8b0[12]),
    .o(al_d6e945fd[12]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e8fb3022 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[7]),
    .c(al_2422b44d[12]),
    .o(al_43cdfb95));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8d903b65 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[7]),
    .c(al_9c80d3c6[12]),
    .o(al_f152e67e[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_c29546d (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_d3f078c4),
    .d(al_43cdfb95),
    .e(al_d6e945fd[12]),
    .f(al_f152e67e[12]),
    .o(al_786f2a14[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_63593b4 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[8]),
    .c(al_5d3f410a[8]),
    .o(al_58fb4752[8]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_fd6a52a (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[8]),
    .c(al_3c07b31a[13]),
    .o(al_9abe6c71));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fe0d8faf (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[8]),
    .c(al_fbcce8b0[13]),
    .o(al_d6e945fd[13]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_3ac68472 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[8]),
    .c(al_2422b44d[13]),
    .o(al_432fdaf9));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1977e7c0 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[8]),
    .c(al_9c80d3c6[13]),
    .o(al_f152e67e[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_cd3a8421 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_9abe6c71),
    .d(al_432fdaf9),
    .e(al_d6e945fd[13]),
    .f(al_f152e67e[13]),
    .o(al_786f2a14[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ed2f3000 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[9]),
    .c(al_5d3f410a[9]),
    .o(al_58fb4752[9]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_423bffc3 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[9]),
    .c(al_3c07b31a[14]),
    .o(al_17aaf618));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2797414b (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[9]),
    .c(al_fbcce8b0[14]),
    .o(al_d6e945fd[14]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_fc1ed3c3 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[9]),
    .c(al_2422b44d[14]),
    .o(al_5d48c7c5));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2247a3e2 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[9]),
    .c(al_9c80d3c6[14]),
    .o(al_f152e67e[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_f5df92b9 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_17aaf618),
    .d(al_5d48c7c5),
    .e(al_d6e945fd[14]),
    .f(al_f152e67e[14]),
    .o(al_786f2a14[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a99e4df1 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[10]),
    .c(al_5d3f410a[10]),
    .o(al_58fb4752[10]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_e80f95fb (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[10]),
    .c(al_3c07b31a[15]),
    .o(al_10938478));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4dc2faf3 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[10]),
    .c(al_fbcce8b0[15]),
    .o(al_d6e945fd[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_4971520c (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[10]),
    .c(al_2422b44d[15]),
    .o(al_73e027c6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_dd27f333 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[10]),
    .c(al_9c80d3c6[15]),
    .o(al_f152e67e[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_966e20c9 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_10938478),
    .d(al_73e027c6),
    .e(al_d6e945fd[15]),
    .f(al_f152e67e[15]),
    .o(al_786f2a14[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8c7b4e85 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[11]),
    .c(al_5d3f410a[11]),
    .o(al_58fb4752[11]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b5d58990 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[11]),
    .c(al_3c07b31a[16]),
    .o(al_87d947b1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6df1082a (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[11]),
    .c(al_fbcce8b0[16]),
    .o(al_d6e945fd[16]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_db2801c2 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[11]),
    .c(al_2422b44d[16]),
    .o(al_5381ba5b));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_232fef7e (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[11]),
    .c(al_9c80d3c6[16]),
    .o(al_f152e67e[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_254634e5 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_87d947b1),
    .d(al_5381ba5b),
    .e(al_d6e945fd[16]),
    .f(al_f152e67e[16]),
    .o(al_786f2a14[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_208325da (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[12]),
    .c(al_5d3f410a[12]),
    .o(al_58fb4752[12]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_57910267 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[12]),
    .c(al_3c07b31a[17]),
    .o(al_4577c722));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_453b6843 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[12]),
    .c(al_fbcce8b0[17]),
    .o(al_d6e945fd[17]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_5644874 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[12]),
    .c(al_2422b44d[17]),
    .o(al_73962c09));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a79a051a (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[12]),
    .c(al_9c80d3c6[17]),
    .o(al_f152e67e[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_67d04835 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_4577c722),
    .d(al_73962c09),
    .e(al_d6e945fd[17]),
    .f(al_f152e67e[17]),
    .o(al_786f2a14[17]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b01fe095 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[3]),
    .c(al_3c07b31a[1]),
    .o(al_52be79ea));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a271933a (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[3]),
    .c(al_fbcce8b0[1]),
    .o(al_d6e945fd[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_5a011779 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[3]),
    .c(al_2422b44d[1]),
    .o(al_ea8a5d3e));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_100ca0a4 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[3]),
    .c(al_9c80d3c6[1]),
    .o(al_f152e67e[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_cfc30b29 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_52be79ea),
    .d(al_ea8a5d3e),
    .e(al_d6e945fd[1]),
    .f(al_f152e67e[1]),
    .o(al_786f2a14[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ad542a37 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[13]),
    .c(al_5d3f410a[13]),
    .o(al_58fb4752[13]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_75fa04b0 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[13]),
    .c(al_3c07b31a[24]),
    .o(al_e1f78661));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8c036c31 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[13]),
    .c(al_fbcce8b0[24]),
    .o(al_d6e945fd[24]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_3fa46135 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[13]),
    .c(al_2422b44d[24]),
    .o(al_16866029));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f1f98e1d (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[13]),
    .c(al_9c80d3c6[24]),
    .o(al_f152e67e[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_77fdcdef (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_e1f78661),
    .d(al_16866029),
    .e(al_d6e945fd[24]),
    .f(al_f152e67e[24]),
    .o(al_786f2a14[24]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_64a739d9 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[14]),
    .c(al_5d3f410a[14]),
    .o(al_58fb4752[14]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f5de6cb1 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[14]),
    .c(al_3c07b31a[25]),
    .o(al_332b9a71));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e6b7a5f2 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[14]),
    .c(al_fbcce8b0[25]),
    .o(al_d6e945fd[25]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c554bb1c (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[14]),
    .c(al_2422b44d[25]),
    .o(al_2a694afc));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ee364f29 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[14]),
    .c(al_9c80d3c6[25]),
    .o(al_f152e67e[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_3a4757b0 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_332b9a71),
    .d(al_2a694afc),
    .e(al_d6e945fd[25]),
    .f(al_f152e67e[25]),
    .o(al_786f2a14[25]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_44979fc7 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[15]),
    .c(al_5d3f410a[15]),
    .o(al_58fb4752[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_4e0cd6f9 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[15]),
    .c(al_3c07b31a[26]),
    .o(al_5b4201dc));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c8fc82ab (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[15]),
    .c(al_fbcce8b0[26]),
    .o(al_d6e945fd[26]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_3cb4c5f (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[15]),
    .c(al_2422b44d[26]),
    .o(al_be2cdb9a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f83be44d (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[15]),
    .c(al_9c80d3c6[26]),
    .o(al_f152e67e[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_5b5bfe87 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_5b4201dc),
    .d(al_be2cdb9a),
    .e(al_d6e945fd[26]),
    .f(al_f152e67e[26]),
    .o(al_786f2a14[26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4a4a77fc (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[16]),
    .c(al_5d3f410a[16]),
    .o(al_58fb4752[16]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1b2cda28 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[16]),
    .c(al_3c07b31a[27]),
    .o(al_398c67e1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_aad867b3 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[16]),
    .c(al_fbcce8b0[27]),
    .o(al_d6e945fd[27]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_dc2ce4c (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[16]),
    .c(al_2422b44d[27]),
    .o(al_a59eb56e));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f09ad4a (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[16]),
    .c(al_9c80d3c6[27]),
    .o(al_f152e67e[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_bdf90c91 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_398c67e1),
    .d(al_a59eb56e),
    .e(al_d6e945fd[27]),
    .f(al_f152e67e[27]),
    .o(al_786f2a14[27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_208fee0 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[17]),
    .c(al_5d3f410a[17]),
    .o(al_58fb4752[17]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_2c22e5dc (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[17]),
    .c(al_3c07b31a[28]),
    .o(al_3ea833b1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_68c2c00d (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[17]),
    .c(al_fbcce8b0[28]),
    .o(al_d6e945fd[28]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c6aeba8f (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[17]),
    .c(al_2422b44d[28]),
    .o(al_dafbe78d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f3c43fca (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[17]),
    .c(al_9c80d3c6[28]),
    .o(al_f152e67e[28]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_def5eb01 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_3ea833b1),
    .d(al_dafbe78d),
    .e(al_d6e945fd[28]),
    .f(al_f152e67e[28]),
    .o(al_786f2a14[28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f46f8326 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[18]),
    .c(al_5d3f410a[18]),
    .o(al_58fb4752[18]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1f7b3134 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[18]),
    .c(al_3c07b31a[29]),
    .o(al_ef43c30e));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_83949279 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[18]),
    .c(al_fbcce8b0[29]),
    .o(al_d6e945fd[29]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_75af9244 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[18]),
    .c(al_2422b44d[29]),
    .o(al_724c627b));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_af5f8817 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[18]),
    .c(al_9c80d3c6[29]),
    .o(al_f152e67e[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_ab89a8e3 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_ef43c30e),
    .d(al_724c627b),
    .e(al_d6e945fd[29]),
    .f(al_f152e67e[29]),
    .o(al_786f2a14[29]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f5c16524 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[4]),
    .c(al_3c07b31a[2]),
    .o(al_1c4e8451));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2c03c1ef (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[4]),
    .c(al_fbcce8b0[2]),
    .o(al_d6e945fd[2]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_89817e03 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[4]),
    .c(al_2422b44d[2]),
    .o(al_a3df3136));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_aadd45fe (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[4]),
    .c(al_9c80d3c6[2]),
    .o(al_f152e67e[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_ed512040 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_1c4e8451),
    .d(al_a3df3136),
    .e(al_d6e945fd[2]),
    .f(al_f152e67e[2]),
    .o(al_786f2a14[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f6363731 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[19]),
    .c(al_5d3f410a[19]),
    .o(al_58fb4752[19]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_2a8f5318 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[19]),
    .c(al_3c07b31a[30]),
    .o(al_8860002c));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3c1d9b6d (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[19]),
    .c(al_fbcce8b0[30]),
    .o(al_d6e945fd[30]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_bd57994 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[19]),
    .c(al_2422b44d[30]),
    .o(al_5ffe271b));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_abb5aea7 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[19]),
    .c(al_9c80d3c6[30]),
    .o(al_f152e67e[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_5a721c53 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_8860002c),
    .d(al_5ffe271b),
    .e(al_d6e945fd[30]),
    .f(al_f152e67e[30]),
    .o(al_786f2a14[30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_45960e3c (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[20]),
    .c(al_5d3f410a[20]),
    .o(al_58fb4752[20]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_2d2d6ba3 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[20]),
    .c(al_3c07b31a[31]),
    .o(al_2f6c7b59));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1fde0b15 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[20]),
    .c(al_fbcce8b0[31]),
    .o(al_d6e945fd[31]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f62f846d (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[20]),
    .c(al_2422b44d[31]),
    .o(al_d7dd86a1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_22a8f5f0 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[20]),
    .c(al_9c80d3c6[31]),
    .o(al_f152e67e[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_eb47bd45 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_2f6c7b59),
    .d(al_d7dd86a1),
    .e(al_d6e945fd[31]),
    .f(al_f152e67e[31]),
    .o(al_786f2a14[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_eabcb5ab (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[21]),
    .c(al_5d3f410a[21]),
    .o(al_58fb4752[21]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_af0c5053 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[21]),
    .c(al_3c07b31a[32]),
    .o(al_22b5c5ea));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7ea98a2b (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[21]),
    .c(al_fbcce8b0[32]),
    .o(al_d6e945fd[32]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_4bc35b76 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[21]),
    .c(al_2422b44d[32]),
    .o(al_d70f37f4));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_750cdc39 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[21]),
    .c(al_9c80d3c6[32]),
    .o(al_f152e67e[32]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_592d51c2 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_22b5c5ea),
    .d(al_d70f37f4),
    .e(al_d6e945fd[32]),
    .f(al_f152e67e[32]),
    .o(al_786f2a14[32]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3c01feca (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[22]),
    .c(al_5d3f410a[22]),
    .o(al_58fb4752[22]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f51a52b6 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[22]),
    .c(al_3c07b31a[33]),
    .o(al_8d2646f7));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e38d1c28 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[22]),
    .c(al_fbcce8b0[33]),
    .o(al_d6e945fd[33]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6e94a241 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[22]),
    .c(al_2422b44d[33]),
    .o(al_3ebdb95a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e0d15c78 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[22]),
    .c(al_9c80d3c6[33]),
    .o(al_f152e67e[33]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_297932a3 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_8d2646f7),
    .d(al_3ebdb95a),
    .e(al_d6e945fd[33]),
    .f(al_f152e67e[33]),
    .o(al_786f2a14[33]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6a719130 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[23]),
    .c(al_5d3f410a[23]),
    .o(al_58fb4752[23]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_d7aca870 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[23]),
    .c(al_3c07b31a[34]),
    .o(al_323b4714));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_af5a02cc (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[23]),
    .c(al_fbcce8b0[34]),
    .o(al_d6e945fd[34]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_b03c18c8 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[23]),
    .c(al_2422b44d[34]),
    .o(al_e4d0aba8));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4548e0d2 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[23]),
    .c(al_9c80d3c6[34]),
    .o(al_f152e67e[34]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_36e49a93 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_323b4714),
    .d(al_e4d0aba8),
    .e(al_d6e945fd[34]),
    .f(al_f152e67e[34]),
    .o(al_786f2a14[34]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c9e58842 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[24]),
    .c(al_5d3f410a[24]),
    .o(al_58fb4752[24]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_35bf74fc (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[24]),
    .c(al_3c07b31a[35]),
    .o(al_12aaa92f));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_adda7984 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[24]),
    .c(al_fbcce8b0[35]),
    .o(al_d6e945fd[35]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_cbe608e5 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[24]),
    .c(al_2422b44d[35]),
    .o(al_7b9f0c1d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fd077897 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[24]),
    .c(al_9c80d3c6[35]),
    .o(al_f152e67e[35]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_a23f09ae (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_12aaa92f),
    .d(al_7b9f0c1d),
    .e(al_d6e945fd[35]),
    .f(al_f152e67e[35]),
    .o(al_786f2a14[35]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6608956a (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[25]),
    .c(al_5d3f410a[25]),
    .o(al_58fb4752[25]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_f6fe8d6c (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[25]),
    .c(al_3c07b31a[36]),
    .o(al_2a4334cc));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_86745908 (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[25]),
    .c(al_fbcce8b0[36]),
    .o(al_d6e945fd[36]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_c101e79a (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[25]),
    .c(al_2422b44d[36]),
    .o(al_3ef4ff5b));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_92de8455 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[25]),
    .c(al_9c80d3c6[36]),
    .o(al_f152e67e[36]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_10c4198a (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_2a4334cc),
    .d(al_3ef4ff5b),
    .e(al_d6e945fd[36]),
    .f(al_f152e67e[36]),
    .o(al_786f2a14[36]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a5334acc (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[26]),
    .c(al_5d3f410a[26]),
    .o(al_58fb4752[26]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_7c4a83c4 (
    .a(al_f001c0eb[0]),
    .b(al_58fb4752[26]),
    .c(al_3c07b31a[37]),
    .o(al_e731c778));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_122d0a1a (
    .a(al_f001c0eb[1]),
    .b(al_58fb4752[26]),
    .c(al_fbcce8b0[37]),
    .o(al_d6e945fd[37]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_6ed6d1a4 (
    .a(al_f001c0eb[2]),
    .b(al_58fb4752[26]),
    .c(al_2422b44d[37]),
    .o(al_542b9ee6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_eb2903a9 (
    .a(al_f001c0eb[3]),
    .b(al_58fb4752[26]),
    .c(al_9c80d3c6[37]),
    .o(al_f152e67e[37]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_d07fa05c (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_e731c778),
    .d(al_542b9ee6),
    .e(al_d6e945fd[37]),
    .f(al_f152e67e[37]),
    .o(al_786f2a14[37]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_494ba8b0 (
    .a(ddr_app_rdy),
    .b(al_65621cdc[0]),
    .c(al_bfd664bf[0]),
    .o(al_88a8db2c[0]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_eda3f42a (
    .a(al_f001c0eb[0]),
    .b(al_88a8db2c[0]),
    .c(al_3c07b31a[44]),
    .o(al_3563cff1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a4a1bea (
    .a(al_f001c0eb[1]),
    .b(al_88a8db2c[0]),
    .c(al_fbcce8b0[44]),
    .o(al_d6e945fd[44]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_8c37ed2b (
    .a(al_f001c0eb[2]),
    .b(al_88a8db2c[0]),
    .c(al_2422b44d[44]),
    .o(al_465c1e37));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8d37d23b (
    .a(al_f001c0eb[3]),
    .b(al_88a8db2c[0]),
    .c(al_9c80d3c6[44]),
    .o(al_f152e67e[44]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_35475810 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_3563cff1),
    .d(al_465c1e37),
    .e(al_d6e945fd[44]),
    .f(al_f152e67e[44]),
    .o(al_786f2a14[44]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3bfa95b8 (
    .a(ddr_app_rdy),
    .b(al_65621cdc[1]),
    .c(al_bfd664bf[1]),
    .o(al_88a8db2c[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_df4bf711 (
    .a(al_f001c0eb[0]),
    .b(al_88a8db2c[1]),
    .c(al_3c07b31a[45]),
    .o(al_bc72c85a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d6c6517a (
    .a(al_f001c0eb[1]),
    .b(al_88a8db2c[1]),
    .c(al_fbcce8b0[45]),
    .o(al_d6e945fd[45]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_a6ec29f7 (
    .a(al_f001c0eb[2]),
    .b(al_88a8db2c[1]),
    .c(al_2422b44d[45]),
    .o(al_4904896d));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_17e9384f (
    .a(al_f001c0eb[3]),
    .b(al_88a8db2c[1]),
    .c(al_9c80d3c6[45]),
    .o(al_f152e67e[45]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_4cfadba1 (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_bc72c85a),
    .d(al_4904896d),
    .e(al_d6e945fd[45]),
    .f(al_f152e67e[45]),
    .o(al_786f2a14[45]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_277bd4ef (
    .a(ddr_app_rdy),
    .b(al_65621cdc[2]),
    .c(al_bfd664bf[2]),
    .o(al_88a8db2c[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9b01243a (
    .a(al_f001c0eb[3]),
    .b(al_88a8db2c[2]),
    .c(al_9c80d3c6[46]),
    .o(al_f152e67e[46]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'habef89cd23670145))
    al_8e54aa9d (
    .a(al_e11b20ed[0]),
    .b(al_e11b20ed[1]),
    .c(al_eb1ff054),
    .d(al_5f8ecffd),
    .e(al_d6e945fd[46]),
    .f(al_f152e67e[46]),
    .o(al_786f2a14[46]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_570d796b (
    .a(al_a1373d93[0]),
    .b(al_1124d2df[1]),
    .o(al_f001c0eb[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ae3b08fc (
    .a(al_a1373d93[0]),
    .b(al_a1373d93[1]),
    .o(al_f001c0eb[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_480b1237 (
    .a(al_a1373d93[0]),
    .b(al_a1373d93[1]),
    .o(al_f001c0eb[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5e1525d3 (
    .a(al_a1373d93[0]),
    .b(al_1124d2df[1]),
    .o(al_f001c0eb[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_1cf446b8 (
    .a(al_f001c0eb[0]),
    .b(al_88a8db2c[2]),
    .c(al_3c07b31a[46]),
    .o(al_eb1ff054));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b447428c (
    .a(al_f001c0eb[1]),
    .b(al_88a8db2c[2]),
    .c(al_fbcce8b0[46]),
    .o(al_d6e945fd[46]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_2a4262dc (
    .a(al_f001c0eb[2]),
    .b(al_88a8db2c[2]),
    .c(al_2422b44d[46]),
    .o(al_5f8ecffd));
  AL_DFF_0 al_e374ba6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cb1ca191),
    .en(1'b1),
    .sr(al_4dd68878),
    .ss(1'b0),
    .q(al_f5b9a4c5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_39894b2f (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[0]),
    .d(al_fea7bbd9[0]),
    .e(al_16b7523e[0]),
    .f(al_f82ace94[0]),
    .o(al_4e72a5eb));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_1b1402b1 (
    .a(al_9d2be50d[0]),
    .b(al_9d2be50d[1]),
    .o(al_382cf878));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_4db5f083 (
    .a(al_41c51f8),
    .b(al_ce2e94ee),
    .c(al_bc5117fe),
    .d(al_8fd7f3b8),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_dc12b1d7));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_54817e9 (
    .a(al_c64ad91c),
    .b(al_5ae0756d),
    .c(al_ef35f7b6[0]),
    .o(al_b59e0dbf));
  AL_MAP_LUT6 #(
    .EQN("(F@~(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'hf0cc55550f33aaaa))
    al_d437b725 (
    .a(al_b59e0dbf),
    .b(al_7eff70ba),
    .c(al_a0f5de0d),
    .d(al_ef35f7b6[0]),
    .e(al_ef35f7b6[1]),
    .f(al_ef35f7b6[34]),
    .o(al_6d82e9d5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_e1821b5e (
    .a(al_b63d0e11),
    .b(al_46d55200),
    .c(al_7e44c8d5),
    .d(al_f7549f58),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_a6bfe69c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_7ce97241 (
    .a(al_2819b010),
    .b(al_98c513dd),
    .c(al_74066232),
    .d(al_f3529ba5),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_a09b37ae));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_2a26166e (
    .a(al_49679814),
    .b(al_c2e0ff4),
    .c(al_bc7b13ca),
    .d(al_7564e3b0),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_6e8781e4));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_388c36ea (
    .a(al_884f3fa8),
    .b(al_91bd4a18),
    .c(al_ef35f7b6[0]),
    .o(al_8a0d8763));
  AL_MAP_LUT6 #(
    .EQN("(F@~(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'hf0cc55550f33aaaa))
    al_6291fd0 (
    .a(al_8a0d8763),
    .b(al_1b5b7fb8),
    .c(al_3f998e21),
    .d(al_ef35f7b6[0]),
    .e(al_ef35f7b6[1]),
    .f(al_ef35f7b6[30]),
    .o(al_afc586c3));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_e44b55c7 (
    .a(al_b169d8ec),
    .b(al_44e6dfe9),
    .c(al_92d8fd60),
    .d(al_7059c89d),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_4c7c6ba3));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_74209d9e (
    .a(al_4e72a5eb),
    .b(al_d149d704),
    .c(al_ef35f7b6[0]),
    .o(al_7040e81f[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_3216a15b (
    .a(al_9c4782d2),
    .b(al_b091346b),
    .c(al_126719a0),
    .d(al_ed48bce4),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_d1e349fb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_4200e746 (
    .a(al_3d92dfa6),
    .b(al_e4f5dc3f),
    .c(al_e8289617),
    .d(al_6b5d2018),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_5fff4931));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_da364cb9 (
    .a(al_13d7dde4),
    .b(al_4c19e182),
    .c(al_ef35f7b6[0]),
    .o(al_ce21c0de));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_957a0ad0 (
    .a(al_ce21c0de),
    .b(al_316deb29),
    .c(al_2115cf8f),
    .d(al_ef35f7b6[0]),
    .e(al_ef35f7b6[1]),
    .f(al_ef35f7b6[31]),
    .o(al_5ea47e0d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_34f743c0 (
    .a(al_4aecdf04),
    .b(al_dcf6b718),
    .c(al_91941257),
    .d(al_47aa4bf9),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_263ba241));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_ed4f8b62 (
    .a(al_2024cd4b),
    .b(al_4e84d779),
    .c(al_df5d8efd),
    .d(al_5758806f),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_50bc0ffd));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_e054e22 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[1]),
    .d(al_fea7bbd9[1]),
    .e(al_16b7523e[1]),
    .f(al_f82ace94[1]),
    .o(al_c307b680));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_92dcbdb7 (
    .a(al_2f7a19ec),
    .b(al_d301de48),
    .c(al_963a39c1),
    .d(al_3f2ddb8a),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_440bddc2));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_c64dbf44 (
    .a(al_c81413d1),
    .b(al_5f6a6401),
    .c(al_ef35f7b6[0]),
    .o(al_bbc46aee));
  AL_MAP_LUT6 #(
    .EQN("(F@(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E))"),
    .INIT(64'h0f33aaaaf0cc5555))
    al_181dd057 (
    .a(al_bbc46aee),
    .b(al_9bbade9e),
    .c(al_3bcdd651),
    .d(al_ef35f7b6[0]),
    .e(al_ef35f7b6[1]),
    .f(al_ef35f7b6[35]),
    .o(al_4ee2ea2f));
  AL_MAP_LUT6 #(
    .EQN("((D@C)*(F@B)*(E@A))"),
    .INIT(64'h0110022004400880))
    al_d2bbfc40 (
    .a(al_4c7c6ba3),
    .b(al_5fff4931),
    .c(al_440bddc2),
    .d(al_ef35f7b6[24]),
    .e(al_ef35f7b6[26]),
    .f(al_ef35f7b6[28]),
    .o(al_932fd4e1));
  AL_MAP_LUT6 #(
    .EQN("(~B*A*(F@D)*(E@C))"),
    .INIT(64'h0002002002002000))
    al_f8f219a3 (
    .a(al_afc586c3),
    .b(al_4ee2ea2f),
    .c(al_a6bfe69c),
    .d(al_50bc0ffd),
    .e(al_ef35f7b6[32]),
    .f(al_ef35f7b6[37]),
    .o(al_eaa2008b));
  AL_MAP_LUT6 #(
    .EQN("((E@C)*(F@B)*(D@A))"),
    .INIT(64'h0102102004084080))
    al_e5b7f0ff (
    .a(al_dc12b1d7),
    .b(al_6e8781e4),
    .c(al_d1e349fb),
    .d(al_ef35f7b6[25]),
    .e(al_ef35f7b6[27]),
    .f(al_ef35f7b6[29]),
    .o(al_2112d3be));
  AL_MAP_LUT6 #(
    .EQN("(~B*A*(F@D)*(E@C))"),
    .INIT(64'h0002002002002000))
    al_92124905 (
    .a(al_6d82e9d5),
    .b(al_5ea47e0d),
    .c(al_a09b37ae),
    .d(al_263ba241),
    .e(al_ef35f7b6[33]),
    .f(al_ef35f7b6[36]),
    .o(al_ceb1b34b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_23ce896e (
    .a(al_5c1c29ee),
    .b(al_9d99a742),
    .c(al_1001936c),
    .d(al_c61f1e9a),
    .e(al_ef35f7b6[0]),
    .f(al_ef35f7b6[1]),
    .o(al_82001be8));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*~B))"),
    .INIT(16'h0405))
    al_d8acb321 (
    .a(al_82001be8),
    .b(al_3e56391),
    .c(al_c088e9dc),
    .d(al_12521532),
    .o(al_1549e910));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_2c9ec636 (
    .a(al_eaa2008b),
    .b(al_ceb1b34b),
    .c(al_932fd4e1),
    .d(al_2112d3be),
    .e(al_1549e910),
    .f(al_382cf878),
    .o(al_d7badb25));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(E*C*B*~A))"),
    .INIT(32'h00bf00ff))
    al_d07b7dae (
    .a(al_c088e9dc),
    .b(al_9d2be50d[0]),
    .c(al_9d2be50d[1]),
    .d(al_9d2be50d[2]),
    .e(al_c360bf4c[3]),
    .o(al_c693d245));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_679c7067 (
    .a(al_c307b680),
    .b(al_d149d704),
    .c(al_ef35f7b6[1]),
    .o(al_7040e81f[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_7b208e69 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[45]),
    .d(al_fea7bbd9[45]),
    .e(al_16b7523e[45]),
    .f(al_f82ace94[45]),
    .o(al_3bbe144d));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_2b845c9 (
    .a(al_3bbe144d),
    .b(al_d149d704),
    .c(al_ef35f7b6[45]),
    .o(al_3242da44));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_eb9f1bb4 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[46]),
    .d(al_fea7bbd9[46]),
    .e(al_16b7523e[46]),
    .f(al_f82ace94[46]),
    .o(al_9c2c924a));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_93ad8f40 (
    .a(al_9c2c924a),
    .b(al_d149d704),
    .c(al_ef35f7b6[46]),
    .o(al_7040e81f[46]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_227a80d4 (
    .a(al_a196b5f4[0]),
    .b(al_a196b5f4[1]),
    .c(al_974136cc[44]),
    .d(al_fea7bbd9[44]),
    .e(al_16b7523e[44]),
    .f(al_f82ace94[44]),
    .o(al_ec32a98f));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_eae2561e (
    .a(init_calib_complete),
    .b(al_90d84dc7[3]),
    .c(al_61f44420),
    .d(ddr_app_rdy),
    .o(al_3e56391));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_8bcecd9 (
    .a(al_ec32a98f),
    .b(al_d149d704),
    .c(al_ef35f7b6[44]),
    .o(al_bc6dea5));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d8db2e85 (
    .a(al_7040e81f[46]),
    .b(al_bc6dea5),
    .o(al_238af9ad));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_fd656049 (
    .a(al_7040e81f[0]),
    .b(al_7040e81f[1]),
    .c(al_63204f4),
    .d(al_6f5534a0),
    .e(al_f1c7f7af),
    .f(al_cf38d855),
    .o(al_43f6f764));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~(~D*~(C*~A))))"),
    .INIT(32'h00233333))
    al_41fe13ed (
    .a(al_d7badb25),
    .b(al_43f6f764),
    .c(al_c693d245),
    .d(al_edebd92e),
    .e(al_d149d704),
    .o(al_8e6a6170));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_89d1c2b9 (
    .a(al_238af9ad),
    .b(al_3242da44),
    .o(al_fc44176c));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_bfd585c9 (
    .a(al_3242da44),
    .b(al_7040e81f[46]),
    .c(al_bc6dea5),
    .d(al_10aff3dd[0]),
    .e(al_10aff3dd[1]),
    .o(al_9609e9f9));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    al_45e18509 (
    .a(al_c088e9dc),
    .b(al_9d2be50d[0]),
    .c(al_9d2be50d[1]),
    .d(al_9d2be50d[2]),
    .o(al_edebd92e));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~(C*~B*A)))"),
    .INIT(32'h00ff0020))
    al_5d1d5f87 (
    .a(al_8e6a6170),
    .b(al_fc44176c),
    .c(al_9609e9f9),
    .d(al_d51c2ed1),
    .e(al_f5b9a4c5),
    .o(al_cb1ca191));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_84ab715 (
    .i(al_a3c26eaf),
    .o(al_8e0772e5));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c445e5ba (
    .i(al_8e0772e5),
    .o(al_b5a5e144));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    al_71651c0b (
    .a(al_60bb426f),
    .b(al_a91e0413[1]),
    .c(al_ee18df00[1]),
    .d(al_ee18df00[0]),
    .o(al_71a56a93[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf6b2d490))
    al_2bd2bf4c (
    .a(al_60bb426f),
    .b(al_a91e0413[1]),
    .c(al_ee18df00[1]),
    .d(al_ee18df00[2]),
    .e(al_ee18df00[0]),
    .o(al_f05e4262[1]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd64b920))
    al_9ff67349 (
    .a(al_60bb426f),
    .b(al_a91e0413[1]),
    .c(al_ee18df00[1]),
    .d(al_ee18df00[2]),
    .e(al_ee18df00[3]),
    .o(al_f05e4262[2]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd64b920))
    al_dfd5d05a (
    .a(al_60bb426f),
    .b(al_a91e0413[1]),
    .c(al_ee18df00[2]),
    .d(al_ee18df00[3]),
    .e(al_ee18df00[4]),
    .o(al_f05e4262[3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hbb20))
    al_bca66adb (
    .a(al_60bb426f),
    .b(al_a91e0413[1]),
    .c(al_ee18df00[3]),
    .d(al_ee18df00[4]),
    .o(al_f05e4262[4]));
  AL_DFF_0 al_6d3f2266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c2672a0d),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a91e0413[0]));
  AL_DFF_0 al_31a1e66e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a91e0413[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a91e0413[1]));
  AL_DFF_0 al_1b148bcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f05e4262[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_ee18df00[4]));
  AL_DFF_1 al_3ed55ad7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71a56a93[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(al_b5a5e144),
    .q(al_ee18df00[0]));
  AL_DFF_0 al_c9901f08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f05e4262[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_ee18df00[1]));
  AL_DFF_0 al_2d29b1f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f05e4262[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_ee18df00[2]));
  AL_DFF_0 al_cda5d34e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f05e4262[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_ee18df00[3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D)"),
    .INIT(16'h0116))
    al_98eb1816 (
    .a(al_c360bf4c[0]),
    .b(al_c360bf4c[1]),
    .c(al_c360bf4c[2]),
    .d(al_c360bf4c[3]),
    .o(al_c2672a0d));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_46a6a3de (
    .a(al_edb1c8b0),
    .b(al_ee18df00[4]),
    .c(al_c360bf4c[1]),
    .o(al_a8be2de9[1]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    al_a4a7a433 (
    .a(al_a8be2de9[1]),
    .b(al_71e16f2b),
    .c(al_ee18df00[4]),
    .d(al_c360bf4c[0]),
    .o(al_43519c87));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_15d64ef0 (
    .a(al_1c8747c7),
    .b(al_ee18df00[4]),
    .c(al_c360bf4c[3]),
    .o(al_a8be2de9[3]));
  AL_MAP_LUT5 #(
    .EQN("~(~B*A*~(~E*~D*C))"),
    .INIT(32'hddddddfd))
    al_e936cbe (
    .a(al_43519c87),
    .b(al_a8be2de9[3]),
    .c(al_15ca36a),
    .d(al_ee18df00[4]),
    .e(al_c360bf4c[2]),
    .o(al_60bb426f));
  AL_MAP_LUT6 #(
    .EQN("(~(~(~F*~D*C)*~B)*~(E*~A))"),
    .INIT(64'h8888cccc88a8ccfc))
    al_9e82aaa0 (
    .a(al_43519c87),
    .b(al_a8be2de9[3]),
    .c(al_15ca36a),
    .d(al_ee18df00[4]),
    .e(al_7f2ef1df),
    .f(al_c360bf4c[2]),
    .o(al_ca609b89));
  AL_MAP_LUT6 #(
    .EQN("(C*~B*A*~(~F*E*D))"),
    .INIT(64'h2020202000202020))
    al_cb489401 (
    .a(al_60bb426f),
    .b(al_ca609b89),
    .c(al_a8be2de9[1]),
    .d(al_71e16f2b),
    .e(al_a92e1411),
    .f(al_c360bf4c[0]),
    .o(al_1a7e2632));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(~C*B)))"),
    .INIT(16'hfbaa))
    al_8abf1228 (
    .a(al_1a7e2632),
    .b(al_60bb426f),
    .c(al_ca609b89),
    .d(al_a92e1411),
    .o(al_d656ab9));
  AL_DFF_0 al_250c614d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d656ab9),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a92e1411));
  AL_MAP_LUT5 #(
    .EQN("(B*A*~(~E*D*C))"),
    .INIT(32'h88880888))
    al_3b2194b4 (
    .a(al_ca609b89),
    .b(al_a8be2de9[3]),
    .c(al_15ca36a),
    .d(al_6748cc6a),
    .e(al_c360bf4c[2]),
    .o(al_618346d9));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    al_3dae64cf (
    .a(al_618346d9),
    .b(al_ca609b89),
    .c(al_6748cc6a),
    .o(al_1e6583f2));
  AL_DFF_0 al_e061722 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1e6583f2),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_6748cc6a));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    al_af19cc8 (
    .a(al_60bb426f),
    .b(al_ca609b89),
    .c(al_7f2ef1df),
    .o(al_93fe255e));
  AL_DFF_0 al_bb50e8b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_93fe255e),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_7f2ef1df));
  AL_DFF_0 al_2855e3a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_176f9515),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c360bf4c[0]));
  AL_DFF_0 al_60f37173 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a7e2632),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c360bf4c[1]));
  AL_DFF_0 al_76b50678 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3bdcd136),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c360bf4c[2]));
  AL_DFF_0 al_49f48857 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_618346d9),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c360bf4c[3]));
  AL_DFF_0 al_b392b9fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_60bb426f),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_1ffff680));
  AL_MAP_LUT6 #(
    .EQN("(~F*C*~A*(~D*~(E)*~(B)+~D*E*~(B)+~(~D)*E*B+~D*E*B))"),
    .INIT(64'h0000000040500010))
    al_fe773c75 (
    .a(al_ca609b89),
    .b(al_a8be2de9[1]),
    .c(al_71e16f2b),
    .d(al_ee18df00[4]),
    .e(al_a92e1411),
    .f(al_c360bf4c[0]),
    .o(al_176f9515));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*~(~E*D*C)))"),
    .INIT(32'h2222a222))
    al_edef6bbb (
    .a(al_ca609b89),
    .b(al_a8be2de9[3]),
    .c(al_15ca36a),
    .d(al_6748cc6a),
    .e(al_c360bf4c[2]),
    .o(al_3bdcd136));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    al_12fb2d87 (
    .a(al_be11f694),
    .b(al_ef9accde),
    .c(al_c58b049c),
    .o(al_9120ce24));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*~(E*~D*C)))"),
    .INIT(32'h22a22222))
    al_f74b3967 (
    .a(al_198de9a1),
    .b(al_a26c7aae[3]),
    .c(al_be11f694),
    .d(al_ef9accde),
    .e(al_c58b049c),
    .o(al_887856fc[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_3953403c (
    .a(al_ef9accde),
    .b(al_5bb559f0),
    .c(al_c9d121b2),
    .o(al_1c402ea2));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_e51e6775 (
    .a(al_ef78cbcb),
    .b(al_1c402ea2),
    .c(al_a70d3eb4),
    .o(al_99fcd329));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_ba64cfb1 (
    .a(al_887856fc[3]),
    .b(al_1c402ea2),
    .o(al_1f4cc6b));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(~A*~(D*~B)))"),
    .INIT(16'h4f5f))
    al_dc2b1 (
    .a(al_887856fc[3]),
    .b(al_ef78cbcb),
    .c(al_1c402ea2),
    .d(al_a70d3eb4),
    .o(al_1846303e));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    al_e4101c6e (
    .a(al_81c227e0[0]),
    .b(al_be11f694),
    .c(al_ef9accde),
    .d(al_c58b049c),
    .o(al_1e3dbb5f));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_df662c77 (
    .a(al_887856fc[0]),
    .b(al_1c402ea2),
    .o(al_c20d9298));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_528a543d (
    .a(al_b4c6b3bd),
    .b(al_1c402ea2),
    .c(al_d50c8b50),
    .o(al_54588780));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(~A*~(D*~B)))"),
    .INIT(16'h4f5f))
    al_a23a256e (
    .a(al_887856fc[0]),
    .b(al_b4c6b3bd),
    .c(al_1c402ea2),
    .d(al_d50c8b50),
    .o(al_a846796e));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*~A)"),
    .INIT(32'h00100000))
    al_6f03da8e (
    .a(al_ef78cbcb),
    .b(al_9120ce24),
    .c(al_f419b7f2),
    .d(al_3f592f2c),
    .e(al_54b33a69),
    .o(al_7ead2bfc[2]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*~A)"),
    .INIT(32'h00100000))
    al_befec5ef (
    .a(al_d51c2ed1),
    .b(al_9120ce24),
    .c(al_f5b9a4c5),
    .d(al_3f592f2c),
    .e(al_54b33a69),
    .o(al_7ead2bfc[3]));
  AL_MAP_LUT6 #(
    .EQN("(~D*~A*~(C*B*~(~F*~E)))"),
    .INIT(64'h0015001500150055))
    al_fe9a0b4f (
    .a(al_1f4cc6b),
    .b(al_1846303e),
    .c(al_a846796e),
    .d(al_99fcd329),
    .e(al_7ead2bfc[2]),
    .f(al_7ead2bfc[3]),
    .o(al_4a7b60f));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*~A)"),
    .INIT(32'h00100000))
    al_2ab84644 (
    .a(al_1e3dbb5f),
    .b(al_9120ce24),
    .c(al_bb796872),
    .d(al_3f592f2c),
    .e(al_54b33a69),
    .o(al_7ead2bfc[0]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*~A)"),
    .INIT(32'h00100000))
    al_713eb2c0 (
    .a(al_b4c6b3bd),
    .b(al_9120ce24),
    .c(al_891497d5),
    .d(al_3f592f2c),
    .e(al_54b33a69),
    .o(al_7ead2bfc[1]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*B*A))"),
    .INIT(16'h070f))
    al_c244a3ee (
    .a(al_1846303e),
    .b(al_a846796e),
    .c(al_54588780),
    .d(al_7ead2bfc[1]),
    .o(al_86879761));
  AL_MAP_LUT6 #(
    .EQN("(~D*~B*~(C*A*~(~F*~E)))"),
    .INIT(64'h0013001300130033))
    al_71183025 (
    .a(al_1846303e),
    .b(al_c20d9298),
    .c(al_a846796e),
    .d(al_54588780),
    .e(al_7ead2bfc[0]),
    .f(al_7ead2bfc[1]),
    .o(al_aed918ac));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~B*~(D*C*A)))"),
    .INIT(32'heccc0000))
    al_6255076f (
    .a(al_1846303e),
    .b(al_c20d9298),
    .c(al_a846796e),
    .d(al_7ead2bfc[0]),
    .e(al_d5d22300),
    .o(al_31deb4f1));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_16306094 (
    .a(al_86879761),
    .b(al_31deb4f1),
    .o(al_bc9b7e1e[1]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(C)*~(D)*~((~E*~B))+A*C*~(D)*~((~E*~B))+A*~(C)*D*~((~E*~B))+~(A)*C*D*~((~E*~B))+A*C*D*~((~E*~B))+~(A)*~(C)*D*(~E*~B)+A*~(C)*D*(~E*~B)+~(A)*C*D*(~E*~B)+A*C*D*(~E*~B))"),
    .INIT(32'hfaaafb88))
    al_b663e6b9 (
    .a(al_bc9b7e1e[1]),
    .b(al_4a7b60f),
    .c(al_aed918ac),
    .d(al_d5d22300),
    .e(al_c30bbc78),
    .o(al_b6f81c2e));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*~(E*~D*C)))"),
    .INIT(32'h22a22222))
    al_af7768ac (
    .a(al_1c1fb07a),
    .b(al_81c227e0[0]),
    .c(al_be11f694),
    .d(al_ef9accde),
    .e(al_c58b049c),
    .o(al_887856fc[0]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    al_feec8971 (
    .a(al_a26c7aae[1]),
    .b(al_be11f694),
    .c(al_ef9accde),
    .d(al_c58b049c),
    .o(al_b4c6b3bd));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    al_267ee063 (
    .a(al_a26c7aae[2]),
    .b(al_be11f694),
    .c(al_ef9accde),
    .d(al_c58b049c),
    .o(al_ef78cbcb));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    al_58602201 (
    .a(al_a26c7aae[3]),
    .b(al_be11f694),
    .c(al_ef9accde),
    .d(al_c58b049c),
    .o(al_d51c2ed1));
  AL_DFF_0 al_dd012eb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6f81c2e),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d5d22300));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a88c44ad (
    .a(al_8704f4a0),
    .b(al_d4979c57),
    .c(al_712d892b),
    .o(al_c8887654));
  AL_DFF_0 al_b8c1a34a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c8887654),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_712d892b));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_bfe9648e (
    .a(al_4a7b60f),
    .b(al_aed918ac),
    .c(al_c30bbc78),
    .o(al_48488f01));
  AL_DFF_0 al_8ec98617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_48488f01),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c30bbc78));
  AL_DFF_0 al_bde6ba94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c4e3d21b),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_81c227e0[0]));
  AL_DFF_0 al_6596bc73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_666055dd),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a26c7aae[1]));
  AL_DFF_0 al_28a089a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69127009),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a26c7aae[2]));
  AL_DFF_0 al_cd79b165 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6a352978),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a26c7aae[3]));
  AL_DFF_0 al_128a8296 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_984f095b[0]),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_aa505777[0]));
  AL_DFF_0 al_c8feefcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_984f095b[1]),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_aa505777[1]));
  AL_DFF_0 al_678ecb19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d53ceeb6[0]),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_1692563a[0]));
  AL_DFF_0 al_fcb8dea1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_24e0f545),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_be11f694));
  AL_MAP_LUT6 #(
    .EQN("(E*~B*~(~D*~C)*~(~F*~A))"),
    .INIT(64'h3330000022200000))
    al_5be0c544 (
    .a(al_4a7b60f),
    .b(al_aed918ac),
    .c(al_86879761),
    .d(al_31deb4f1),
    .e(al_7ead2bfc[0]),
    .f(al_c30bbc78),
    .o(al_ab3d1147));
  AL_MAP_LUT5 #(
    .EQN("(D*~C*~B*~(~E*~A))"),
    .INIT(32'h03000200))
    al_8604807d (
    .a(al_4a7b60f),
    .b(al_86879761),
    .c(al_31deb4f1),
    .d(al_7ead2bfc[1]),
    .e(al_c30bbc78),
    .o(al_a2d1acac));
  AL_MAP_LUT6 #(
    .EQN("~(~C*~B*~(A*(E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)))"),
    .INIT(64'hfefefefcfcfefcfc))
    al_cba7eb38 (
    .a(al_8704f4a0),
    .b(al_ab3d1147),
    .c(al_a2d1acac),
    .d(al_d4979c57),
    .e(al_7ead2bfc[2]),
    .f(al_7ead2bfc[3]),
    .o(al_9d55a7e5));
  AL_DFF_0 al_26905d27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9d55a7e5),
    .en(al_f88e71cf),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_ef9accde));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    al_d48fb970 (
    .a(al_1846303e),
    .b(al_a846796e),
    .o(al_24e0f545));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h080d080cddddcccc))
    al_3ff8cbe5 (
    .a(al_24e0f545),
    .b(al_1f4cc6b),
    .c(al_99fcd329),
    .d(al_7ead2bfc[2]),
    .e(al_7ead2bfc[3]),
    .f(al_712d892b),
    .o(al_d4979c57));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    al_aee3f219 (
    .a(al_4a7b60f),
    .b(al_aed918ac),
    .c(al_c30bbc78),
    .o(al_8704f4a0));
  AL_MAP_LUT6 #(
    .EQN("(E*~B*~(~D*~C)*~(~F*~A))"),
    .INIT(64'h3330000022200000))
    al_23f20a20 (
    .a(al_4a7b60f),
    .b(al_aed918ac),
    .c(al_86879761),
    .d(al_31deb4f1),
    .e(al_31adf876[0]),
    .f(al_c30bbc78),
    .o(al_72131b80));
  AL_MAP_LUT5 #(
    .EQN("(D*~C*~B*~(~E*~A))"),
    .INIT(32'h03000200))
    al_45949f24 (
    .a(al_4a7b60f),
    .b(al_86879761),
    .c(al_31deb4f1),
    .d(al_fd46e088[0]),
    .e(al_c30bbc78),
    .o(al_f436c091));
  AL_MAP_LUT6 #(
    .EQN("~(~C*~B*~(A*(E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)))"),
    .INIT(64'hfefefefcfcfefcfc))
    al_c8a7d478 (
    .a(al_8704f4a0),
    .b(al_72131b80),
    .c(al_f436c091),
    .d(al_d4979c57),
    .e(al_aaf3456[0]),
    .f(al_4ed70d21[0]),
    .o(al_984f095b[0]));
  AL_MAP_LUT6 #(
    .EQN("(E*~B*~(~D*~C)*~(~F*~A))"),
    .INIT(64'h3330000022200000))
    al_c376f3e2 (
    .a(al_4a7b60f),
    .b(al_aed918ac),
    .c(al_86879761),
    .d(al_31deb4f1),
    .e(al_31adf876[1]),
    .f(al_c30bbc78),
    .o(al_4c923ed));
  AL_MAP_LUT5 #(
    .EQN("(D*~C*~B*~(~E*~A))"),
    .INIT(32'h03000200))
    al_b493bb51 (
    .a(al_4a7b60f),
    .b(al_86879761),
    .c(al_31deb4f1),
    .d(al_fd46e088[1]),
    .e(al_c30bbc78),
    .o(al_becbe1a2));
  AL_MAP_LUT6 #(
    .EQN("~(~C*~B*~(A*(E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)))"),
    .INIT(64'hfefefefcfcfefcfc))
    al_fa5c5947 (
    .a(al_8704f4a0),
    .b(al_4c923ed),
    .c(al_becbe1a2),
    .d(al_d4979c57),
    .e(al_aaf3456[1]),
    .f(al_4ed70d21[1]),
    .o(al_984f095b[1]));
  AL_MAP_LUT6 #(
    .EQN("(E*~B*~(~D*~C)*~(~F*~A))"),
    .INIT(64'h3330000022200000))
    al_88a46469 (
    .a(al_4a7b60f),
    .b(al_aed918ac),
    .c(al_86879761),
    .d(al_31deb4f1),
    .e(al_d76fa964[0]),
    .f(al_c30bbc78),
    .o(al_adcb2e1b));
  AL_MAP_LUT5 #(
    .EQN("(D*~C*~B*~(~E*~A))"),
    .INIT(32'h03000200))
    al_8774acea (
    .a(al_4a7b60f),
    .b(al_86879761),
    .c(al_31deb4f1),
    .d(al_d76fa964[2]),
    .e(al_c30bbc78),
    .o(al_43250e7c));
  AL_MAP_LUT6 #(
    .EQN("~(~C*~B*~(A*(E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)))"),
    .INIT(64'hfefefefcfcfefcfc))
    al_3315e838 (
    .a(al_8704f4a0),
    .b(al_adcb2e1b),
    .c(al_43250e7c),
    .d(al_d4979c57),
    .e(al_d76fa964[4]),
    .f(al_d76fa964[6]),
    .o(al_d53ceeb6[0]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*~B))"),
    .INIT(16'h0504))
    al_60934d8b (
    .a(al_bc9b7e1e[1]),
    .b(al_4a7b60f),
    .c(al_aed918ac),
    .d(al_c30bbc78),
    .o(al_c4e3d21b));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    al_9d9def8d (
    .a(al_bc9b7e1e[1]),
    .b(al_4a7b60f),
    .c(al_c30bbc78),
    .o(al_666055dd));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_f64156dd (
    .a(al_8704f4a0),
    .b(al_d4979c57),
    .o(al_69127009));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_fc2f8e28 (
    .a(al_8704f4a0),
    .b(al_d4979c57),
    .o(al_6a352978));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_ff86c7fe (
    .a(al_b15eb135),
    .b(al_7af754c1),
    .o(al_c8a2915b));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_41ea3c6f (
    .a(al_9d5bb698),
    .b(al_18e5c731),
    .o(al_570aaefb));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_13b93829 (
    .a(al_10ef1903),
    .b(al_a738798f),
    .o(al_3589ff80));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_594a9c18 (
    .a(al_1abc6e62),
    .b(al_b01ab869),
    .o(al_1aea9b48));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_df25031e (
    .a(al_e395c44e),
    .b(al_a135e827),
    .o(al_4483f4ea));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_22eab3e5 (
    .a(al_caa664ee),
    .b(al_c92d59d9),
    .o(al_9af29299));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_3294aac (
    .a(al_332c02d0),
    .b(al_7a253edf),
    .o(al_af82789));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_228073cd (
    .a(al_781760a2),
    .b(al_13a574fa),
    .o(al_37c023d));
  AL_DFF_0 al_7ff74b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_30565995),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7077f69));
  AL_DFF_0 al_2d3aea39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b71ef602),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d5bb698));
  AL_DFF_0 al_7ccce9f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0a7db18),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_432e33d4));
  AL_DFF_0 al_1e3c2e1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_89d8cddf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_10ef1903));
  AL_DFF_0 al_a8781214 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2242adc3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eaad117a));
  AL_DFF_0 al_5628e47f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aead4311),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1abc6e62));
  AL_DFF_0 al_1da680b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_beed7bdd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c473b6a4));
  AL_DFF_0 al_d51fbd85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fe8a405),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e395c44e));
  AL_DFF_0 al_6e4cd33c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c032a2f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8454367));
  AL_DFF_0 al_e781c91f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a53fdc6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_caa664ee));
  AL_DFF_0 al_96a6de20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c330002d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fd0c8ec3));
  AL_DFF_0 al_659e993c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0693577),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_332c02d0));
  AL_DFF_0 al_27fd4f7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_76e6275e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a8b491ea));
  AL_DFF_0 al_f6375494 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fb080638),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_781760a2));
  AL_DFF_0 al_868e85ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d17319e5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1c83794e));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_cb6ec46b (
    .a(al_8ed48b41[1]),
    .b(al_8941a5fb[1]),
    .c(al_ef35f7b6[1]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_18e4b32e));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_47a200e3 (
    .a(al_18e4b32e),
    .b(al_b93da8d5[1]),
    .c(al_c360bf4c[0]),
    .o(al_96d05ba4));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_46684d51 (
    .a(al_8ed48b41[2]),
    .b(al_8941a5fb[2]),
    .c(al_ef35f7b6[2]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_12c2377a));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_a20f4396 (
    .a(al_12c2377a),
    .b(al_b93da8d5[2]),
    .c(al_c360bf4c[0]),
    .o(al_ed3799e7));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fd2f698a (
    .a(al_ed3799e7),
    .b(al_1ffff680),
    .o(al_779bd70c[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_2fef173d (
    .a(al_8ed48b41[0]),
    .b(al_8941a5fb[0]),
    .c(al_ef35f7b6[0]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_f42e5022));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_e1fe1e2e (
    .a(al_f42e5022),
    .b(al_b93da8d5[0]),
    .c(al_c360bf4c[0]),
    .o(al_837d8da3));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_7e6048f0 (
    .a(al_b5a5e144),
    .b(al_a8b491ea),
    .c(al_781760a2),
    .o(al_76e6275e));
  AL_MAP_LUT6 #(
    .EQN("(~D*~(~(F*E)*~(~C*~B*A)))"),
    .INIT(64'h00ff000200020002))
    al_9de13e88 (
    .a(al_779bd70c[2]),
    .b(al_96d05ba4),
    .c(al_837d8da3),
    .d(al_b5a5e144),
    .e(al_a8b491ea),
    .f(al_781760a2),
    .o(al_fb080638));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_64de2d63 (
    .a(al_b5a5e144),
    .b(al_8454367),
    .c(al_caa664ee),
    .o(al_5c032a2f));
  AL_MAP_LUT6 #(
    .EQN("(~D*~(~(F*E)*~(~C*B*A)))"),
    .INIT(64'h00ff000800080008))
    al_8696c09b (
    .a(al_779bd70c[2]),
    .b(al_96d05ba4),
    .c(al_837d8da3),
    .d(al_b5a5e144),
    .e(al_8454367),
    .f(al_caa664ee),
    .o(al_1a53fdc6));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_7e9b199c (
    .a(al_b5a5e144),
    .b(al_f7077f69),
    .c(al_9d5bb698),
    .o(al_30565995));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_a693e52a (
    .a(al_ed3799e7),
    .b(al_b5a5e144),
    .c(al_1ffff680),
    .o(al_b6bef94));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(~C*B*A))"),
    .INIT(64'h08ff080808080808))
    al_840cdd7c (
    .a(al_b6bef94),
    .b(al_96d05ba4),
    .c(al_837d8da3),
    .d(al_b5a5e144),
    .e(al_f7077f69),
    .f(al_9d5bb698),
    .o(al_b71ef602));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_96fa30f6 (
    .a(al_b5a5e144),
    .b(al_eaad117a),
    .c(al_1abc6e62),
    .o(al_2242adc3));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(~C*~B*A))"),
    .INIT(64'h02ff020202020202))
    al_c8d82861 (
    .a(al_b6bef94),
    .b(al_96d05ba4),
    .c(al_837d8da3),
    .d(al_b5a5e144),
    .e(al_eaad117a),
    .f(al_1abc6e62),
    .o(al_aead4311));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_65f82dbb (
    .a(al_b5a5e144),
    .b(al_1c83794e),
    .c(al_b15eb135),
    .o(al_d17319e5));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(C*B*A))"),
    .INIT(64'h80ff808080808080))
    al_fd5f49b5 (
    .a(al_b6bef94),
    .b(al_96d05ba4),
    .c(al_837d8da3),
    .d(al_b5a5e144),
    .e(al_1c83794e),
    .f(al_b15eb135),
    .o(al_96a05b));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_c68a670a (
    .a(al_b5a5e144),
    .b(al_432e33d4),
    .c(al_10ef1903),
    .o(al_c0a7db18));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(C*~B*A))"),
    .INIT(64'h20ff202020202020))
    al_46670b7e (
    .a(al_b6bef94),
    .b(al_96d05ba4),
    .c(al_837d8da3),
    .d(al_b5a5e144),
    .e(al_432e33d4),
    .f(al_10ef1903),
    .o(al_89d8cddf));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_e961c6ac (
    .a(al_b5a5e144),
    .b(al_c473b6a4),
    .c(al_e395c44e),
    .o(al_beed7bdd));
  AL_MAP_LUT6 #(
    .EQN("(~D*~(~(F*E)*~(C*B*A)))"),
    .INIT(64'h00ff008000800080))
    al_dd2b7a30 (
    .a(al_779bd70c[2]),
    .b(al_96d05ba4),
    .c(al_837d8da3),
    .d(al_b5a5e144),
    .e(al_c473b6a4),
    .f(al_e395c44e),
    .o(al_fe8a405));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_fbf0f262 (
    .a(al_b5a5e144),
    .b(al_fd0c8ec3),
    .c(al_332c02d0),
    .o(al_c330002d));
  AL_MAP_LUT6 #(
    .EQN("(~D*~(~(F*E)*~(C*~B*A)))"),
    .INIT(64'h00ff002000200020))
    al_782b96f4 (
    .a(al_779bd70c[2]),
    .b(al_96d05ba4),
    .c(al_837d8da3),
    .d(al_b5a5e144),
    .e(al_fd0c8ec3),
    .f(al_332c02d0),
    .o(al_c0693577));
  AL_DFF_0 al_4c7eda0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_96a05b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b15eb135));
  AL_DFF_0 al_280a69a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4e6ba179),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a868c71));
  AL_DFF_0 al_71a60e36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_237c733d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18e5c731));
  AL_DFF_0 al_9c69b339 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7d5a8c76),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9650ab3a));
  AL_DFF_0 al_ab32ad26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9b32a85e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a738798f));
  AL_DFF_0 al_61296e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2374b47d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_72b1cb56));
  AL_DFF_0 al_4b1558e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7e2e3620),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b01ab869));
  AL_DFF_0 al_af31e108 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8dc1b606),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9ad2b6c));
  AL_DFF_0 al_ea345c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_35f3cf28),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a135e827));
  AL_DFF_0 al_7711a652 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bfe50c52),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7fa83c38));
  AL_DFF_0 al_b6dd52a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f149b540),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c92d59d9));
  AL_DFF_0 al_d4253746 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_53cd58ac),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8194720));
  AL_DFF_0 al_f94f3209 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b3e9d06c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7a253edf));
  AL_DFF_0 al_24991f9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c84ffce0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_231ef4df));
  AL_DFF_0 al_d4a9b97d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c5d5a3f6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13a574fa));
  AL_DFF_0 al_666ce832 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fb9a605b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_99ca5e59));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_254d4380 (
    .a(al_b5a5e144),
    .b(al_231ef4df),
    .c(al_13a574fa),
    .o(al_c84ffce0));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_bc1f821e (
    .a(al_fd46e088[0]),
    .b(al_aaf3456[0]),
    .c(al_4ed70d21[0]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_6b991e1c));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_732cc16e (
    .a(al_6b991e1c),
    .b(al_31adf876[0]),
    .c(al_81c227e0[0]),
    .o(al_d46ec896));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_75d5eabd (
    .a(al_fd46e088[1]),
    .b(al_aaf3456[1]),
    .c(al_4ed70d21[1]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_5dd540e5));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_1a024d70 (
    .a(al_5dd540e5),
    .b(al_31adf876[1]),
    .c(al_81c227e0[0]),
    .o(al_79f445c4));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_a6f46dfb (
    .a(al_d76fa964[2]),
    .b(al_d76fa964[4]),
    .c(al_d76fa964[6]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_57b41659));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_23ebf6c2 (
    .a(al_57b41659),
    .b(al_d76fa964[0]),
    .c(al_81c227e0[0]),
    .o(al_2d6bf5be));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_4622fdf4 (
    .a(al_2d6bf5be),
    .b(al_b5a5e144),
    .c(al_ef9accde),
    .o(al_842732c2));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(~C*~B*A))"),
    .INIT(64'h02ff020202020202))
    al_ec5f7f6a (
    .a(al_842732c2),
    .b(al_d46ec896),
    .c(al_79f445c4),
    .d(al_b5a5e144),
    .e(al_231ef4df),
    .f(al_13a574fa),
    .o(al_c5d5a3f6));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_6b988a06 (
    .a(al_b5a5e144),
    .b(al_72b1cb56),
    .c(al_b01ab869),
    .o(al_2374b47d));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_dcc9c08d (
    .a(al_2d6bf5be),
    .b(al_b5a5e144),
    .c(al_ef9accde),
    .o(al_b3d60ef7));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(~C*~B*A))"),
    .INIT(64'h02ff020202020202))
    al_b297109d (
    .a(al_b3d60ef7),
    .b(al_d46ec896),
    .c(al_79f445c4),
    .d(al_b5a5e144),
    .e(al_72b1cb56),
    .f(al_b01ab869),
    .o(al_7e2e3620));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_5a5febcb (
    .a(al_b5a5e144),
    .b(al_9650ab3a),
    .c(al_a738798f),
    .o(al_7d5a8c76));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(~C*B*A))"),
    .INIT(64'h08ff080808080808))
    al_1c2136bc (
    .a(al_b3d60ef7),
    .b(al_d46ec896),
    .c(al_79f445c4),
    .d(al_b5a5e144),
    .e(al_9650ab3a),
    .f(al_a738798f),
    .o(al_9b32a85e));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_c7363450 (
    .a(al_b5a5e144),
    .b(al_8194720),
    .c(al_7a253edf),
    .o(al_53cd58ac));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(~C*B*A))"),
    .INIT(64'h08ff080808080808))
    al_d57912a3 (
    .a(al_842732c2),
    .b(al_d46ec896),
    .c(al_79f445c4),
    .d(al_b5a5e144),
    .e(al_8194720),
    .f(al_7a253edf),
    .o(al_b3e9d06c));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_a47312df (
    .a(al_b5a5e144),
    .b(al_99ca5e59),
    .c(al_7af754c1),
    .o(al_fb9a605b));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(C*B*A))"),
    .INIT(64'h80ff808080808080))
    al_b46383fa (
    .a(al_b3d60ef7),
    .b(al_d46ec896),
    .c(al_79f445c4),
    .d(al_b5a5e144),
    .e(al_99ca5e59),
    .f(al_7af754c1),
    .o(al_db7ff57e));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_28547a3b (
    .a(al_b5a5e144),
    .b(al_3a868c71),
    .c(al_18e5c731),
    .o(al_4e6ba179));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(C*~B*A))"),
    .INIT(64'h20ff202020202020))
    al_50ef65aa (
    .a(al_b3d60ef7),
    .b(al_d46ec896),
    .c(al_79f445c4),
    .d(al_b5a5e144),
    .e(al_3a868c71),
    .f(al_18e5c731),
    .o(al_237c733d));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_45e5d4cb (
    .a(al_b5a5e144),
    .b(al_a9ad2b6c),
    .c(al_a135e827),
    .o(al_8dc1b606));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(C*B*A))"),
    .INIT(64'h80ff808080808080))
    al_dbcf343f (
    .a(al_842732c2),
    .b(al_d46ec896),
    .c(al_79f445c4),
    .d(al_b5a5e144),
    .e(al_a9ad2b6c),
    .f(al_a135e827),
    .o(al_35f3cf28));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_df219ff0 (
    .a(al_b5a5e144),
    .b(al_7fa83c38),
    .c(al_c92d59d9),
    .o(al_bfe50c52));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~D)*~(C*~B*A))"),
    .INIT(64'h20ff202020202020))
    al_3380a869 (
    .a(al_842732c2),
    .b(al_d46ec896),
    .c(al_79f445c4),
    .d(al_b5a5e144),
    .e(al_7fa83c38),
    .f(al_c92d59d9),
    .o(al_f149b540));
  AL_DFF_0 al_9f769d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_db7ff57e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af754c1));
  AL_DFF_0 al_1fa6deab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c8a2915b),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_fb5f08ff));
  AL_DFF_0 al_9d508437 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_570aaefb),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_90254f7));
  AL_DFF_0 al_f6e0139c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3589ff80),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_b9ff4892));
  AL_DFF_0 al_b37069be (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1aea9b48),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_63860ff5));
  AL_DFF_0 al_f780361b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4483f4ea),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_15578244));
  AL_DFF_0 al_561b38d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9af29299),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_21e21c));
  AL_DFF_0 al_88fcbaee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_af82789),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_9602e904));
  AL_DFF_0 al_442e2c42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_37c023d),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_6d6f00e5));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_b8d34620 (
    .a(al_b5a5e144),
    .o(al_9388375e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_38cce20a (
    .a(al_53bb123b[6]),
    .b(al_53bb123b[7]),
    .c(al_15578244),
    .d(al_21e21c),
    .e(al_9602e904),
    .f(al_6d6f00e5),
    .o(al_c9eb9f8c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_871b78ec (
    .a(al_53bb123b[0]),
    .b(al_53bb123b[1]),
    .c(al_15578244),
    .d(al_21e21c),
    .e(al_9602e904),
    .f(al_6d6f00e5),
    .o(al_2cd04711));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_4cbf018a (
    .a(al_53bb123b[0]),
    .b(al_53bb123b[1]),
    .c(al_fb5f08ff),
    .d(al_90254f7),
    .e(al_b9ff4892),
    .f(al_63860ff5),
    .o(al_b14bdbb3));
  AL_MAP_LUT5 #(
    .EQN("(~E*C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(32'h000050c0))
    al_4da99bbf (
    .a(al_2cd04711),
    .b(al_b14bdbb3),
    .c(al_c56a3e50),
    .d(al_cbeafa67[0]),
    .e(al_90a0fe97[0]),
    .o(al_f01dcc55));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_b21c572 (
    .a(al_53bb123b[2]),
    .b(al_53bb123b[3]),
    .c(al_15578244),
    .d(al_21e21c),
    .e(al_9602e904),
    .f(al_6d6f00e5),
    .o(al_f13534df));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_2afd3575 (
    .a(al_53bb123b[2]),
    .b(al_53bb123b[3]),
    .c(al_fb5f08ff),
    .d(al_90254f7),
    .e(al_b9ff4892),
    .f(al_63860ff5),
    .o(al_9fccc935));
  AL_MAP_LUT5 #(
    .EQN("(~E*C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(32'h000050c0))
    al_4197675a (
    .a(al_f13534df),
    .b(al_9fccc935),
    .c(al_ef9d2d1b),
    .d(al_cbeafa67[2]),
    .e(al_8932a489),
    .o(al_187c11ca[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_ed0ad0af (
    .a(al_f01dcc55),
    .b(al_187c11ca[1]),
    .o(al_c48ef761));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(~C*~A))"),
    .INIT(8'hcd))
    al_b72d712e (
    .a(al_6f337ab4),
    .b(al_c48ef761),
    .c(al_385080cf),
    .o(al_9e404664));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    al_a836959d (
    .a(al_f01dcc55),
    .b(al_187c11ca[1]),
    .c(al_80f00b),
    .o(al_437ca69f[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bf17d4c0 (
    .a(al_9e404664),
    .b(al_437ca69f[1]),
    .c(al_80f00b),
    .o(al_484d3915));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_1312afd3 (
    .a(al_53bb123b[6]),
    .b(al_53bb123b[7]),
    .c(al_fb5f08ff),
    .d(al_90254f7),
    .e(al_b9ff4892),
    .f(al_63860ff5),
    .o(al_ccd9a7ea));
  AL_MAP_LUT5 #(
    .EQN("(~E*C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(32'h000050c0))
    al_3992df6 (
    .a(al_c9eb9f8c),
    .b(al_ccd9a7ea),
    .c(al_dd965664),
    .d(al_cbeafa67[6]),
    .e(al_4c58e022),
    .o(al_187c11ca[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_27153a37 (
    .a(al_53bb123b[4]),
    .b(al_53bb123b[5]),
    .c(al_15578244),
    .d(al_21e21c),
    .e(al_9602e904),
    .f(al_6d6f00e5),
    .o(al_8c8e8f6a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_610ef8ad (
    .a(al_53bb123b[4]),
    .b(al_53bb123b[5]),
    .c(al_fb5f08ff),
    .d(al_90254f7),
    .e(al_b9ff4892),
    .f(al_63860ff5),
    .o(al_b905b88f));
  AL_MAP_LUT5 #(
    .EQN("(~E*C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(32'h000050c0))
    al_71cca5bd (
    .a(al_8c8e8f6a),
    .b(al_b905b88f),
    .c(al_4135f4fc),
    .d(al_cbeafa67[4]),
    .e(al_165f2734),
    .o(al_ab817290));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_a30fa744 (
    .a(al_187c11ca[3]),
    .b(al_ab817290),
    .o(al_6f337ab4));
  AL_DFF_0 al_9bf2eefd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_484d3915),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_80f00b));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    al_d51065fa (
    .a(al_187c11ca[3]),
    .b(al_ab817290),
    .c(al_198bf41a),
    .o(al_ac2fd07f));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_30287dc1 (
    .a(al_c48ef761),
    .b(al_385080cf),
    .o(al_e7ffa4ec));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfe44))
    al_b29c4107 (
    .a(al_e7ffa4ec),
    .b(al_ac2fd07f),
    .c(al_6f337ab4),
    .d(al_198bf41a),
    .o(al_d39ce0c));
  AL_DFF_0 al_8d72b58f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d39ce0c),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_198bf41a));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_f610c6a1 (
    .a(al_6f337ab4),
    .b(al_c48ef761),
    .c(al_385080cf),
    .o(al_b71b7f68));
  AL_DFF_0 al_fce474d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b71b7f68),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_385080cf));
  AL_DFF_0 al_ea8db818 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fbec08cf),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_90a0fe97[0]));
  AL_DFF_0 al_501ee8b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d3598a31),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_8932a489));
  AL_DFF_0 al_2979bd28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bf3d0760),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_165f2734));
  AL_DFF_0 al_e56f55bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8211c6dd),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_4c58e022));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_8c127d17 (
    .a(al_9e404664),
    .b(al_437ca69f[1]),
    .c(al_f01dcc55),
    .o(al_fbec08cf));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fefd2534 (
    .a(al_9e404664),
    .b(al_437ca69f[1]),
    .o(al_d3598a31));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_88ca6f64 (
    .a(al_e7ffa4ec),
    .b(al_ac2fd07f),
    .c(al_6f337ab4),
    .o(al_bf3d0760));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f37b264f (
    .a(al_e7ffa4ec),
    .b(al_ac2fd07f),
    .o(al_8211c6dd));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_506a9b42 (
    .a(al_8ed48b41[24]),
    .b(al_8941a5fb[24]),
    .c(al_ef35f7b6[24]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_a1fbbbd1));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_cb0a31d7 (
    .a(al_a1fbbbd1),
    .b(al_b93da8d5[24]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_eb9aa630[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_ae6a16aa (
    .a(al_46b8ac3c),
    .b(al_4ba8484b),
    .c(al_4f7a36e8),
    .o(al_eb9aa630[6]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_cd0817d2 (
    .a(al_8ed48b41[34]),
    .b(al_8941a5fb[34]),
    .c(al_ef35f7b6[34]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_58de2ea4));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_cfcb6424 (
    .a(al_58de2ea4),
    .b(al_b93da8d5[34]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_3c0a4ef0[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_592ff90b (
    .a(al_8ed48b41[35]),
    .b(al_8941a5fb[35]),
    .c(al_ef35f7b6[35]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_db15dba5));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_13e048c5 (
    .a(al_db15dba5),
    .b(al_b93da8d5[35]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_ecc8e317[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_930b3851 (
    .a(al_8ed48b41[36]),
    .b(al_8941a5fb[36]),
    .c(al_ef35f7b6[36]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_db39a0bd));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_aa60d876 (
    .a(al_db39a0bd),
    .b(al_b93da8d5[36]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_c8b553c9[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_a811ffd7 (
    .a(al_8ed48b41[37]),
    .b(al_8941a5fb[37]),
    .c(al_ef35f7b6[37]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_c3565be1));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_cd430143 (
    .a(al_c3565be1),
    .b(al_b93da8d5[37]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_92812db2[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_221bfd56 (
    .a(al_8ed48b41[25]),
    .b(al_8941a5fb[25]),
    .c(al_ef35f7b6[25]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_6f81b627));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_948673c4 (
    .a(al_6f81b627),
    .b(al_b93da8d5[25]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_534b111d[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_e2564288 (
    .a(al_8ed48b41[26]),
    .b(al_8941a5fb[26]),
    .c(al_ef35f7b6[26]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_76bac341));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_5807d854 (
    .a(al_76bac341),
    .b(al_b93da8d5[26]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_39691102[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_8458f6f2 (
    .a(al_8ed48b41[27]),
    .b(al_8941a5fb[27]),
    .c(al_ef35f7b6[27]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_588f198a));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_fad04247 (
    .a(al_588f198a),
    .b(al_b93da8d5[27]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_304bc4cf[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_fbdefdae (
    .a(al_8ed48b41[28]),
    .b(al_8941a5fb[28]),
    .c(al_ef35f7b6[28]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_9ac35c50));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_525ed3bf (
    .a(al_9ac35c50),
    .b(al_b93da8d5[28]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_421a630e[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_6e5dc3ae (
    .a(al_8ed48b41[29]),
    .b(al_8941a5fb[29]),
    .c(al_ef35f7b6[29]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_5606bbf4));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_6a36c3f7 (
    .a(al_5606bbf4),
    .b(al_b93da8d5[29]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_2cee9b7b[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_81dc5d81 (
    .a(al_8ed48b41[30]),
    .b(al_8941a5fb[30]),
    .c(al_ef35f7b6[30]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_c993dae4));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_1a72bb61 (
    .a(al_c993dae4),
    .b(al_b93da8d5[30]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_2f77b9ea[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_d47fccbf (
    .a(al_8ed48b41[31]),
    .b(al_8941a5fb[31]),
    .c(al_ef35f7b6[31]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_a06bb9a1));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_a4ee5526 (
    .a(al_a06bb9a1),
    .b(al_b93da8d5[31]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_b7a66cc8[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_a0f25feb (
    .a(al_8ed48b41[32]),
    .b(al_8941a5fb[32]),
    .c(al_ef35f7b6[32]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_4b03c837));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_1b4b69cc (
    .a(al_4b03c837),
    .b(al_b93da8d5[32]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_bce3182d[2]));
  AL_MAP_LUT6 #(
    .EQN("~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'h5533550f553355ff))
    al_79116cc6 (
    .a(al_8ed48b41[33]),
    .b(al_8941a5fb[33]),
    .c(al_ef35f7b6[33]),
    .d(al_c360bf4c[1]),
    .e(al_c360bf4c[2]),
    .f(al_c360bf4c[3]),
    .o(al_f8e44d17));
  AL_MAP_LUT4 #(
    .EQN("(D*(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'hc500))
    al_2c4c8081 (
    .a(al_f8e44d17),
    .b(al_b93da8d5[33]),
    .c(al_c360bf4c[0]),
    .d(al_1ffff680),
    .o(al_636a0d93[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_aed89232 (
    .a(al_a4f25695),
    .b(al_aa505777[0]),
    .o(al_e3639d7e[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f440dc93 (
    .a(al_837d8da3),
    .b(al_1ffff680),
    .o(al_e3639d7e[2]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_45c3c46b (
    .a(al_53bb123b[2]),
    .b(al_53bb123b[4]),
    .c(al_53bb123b[6]),
    .d(al_8932a489),
    .e(al_165f2734),
    .f(al_4c58e022),
    .o(al_a4894768));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_43ec54bc (
    .a(al_a4894768),
    .b(al_53bb123b[0]),
    .c(al_90a0fe97[0]),
    .o(al_e3639d7e[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c9c66c80 (
    .a(al_a4f25695),
    .b(al_aa505777[1]),
    .o(al_18fbbb0f[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_8440aa9f (
    .a(al_96d05ba4),
    .b(al_1ffff680),
    .o(al_18fbbb0f[2]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_c638375 (
    .a(al_53bb123b[3]),
    .b(al_53bb123b[5]),
    .c(al_53bb123b[7]),
    .d(al_8932a489),
    .e(al_165f2734),
    .f(al_4c58e022),
    .o(al_6a408c69));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6614a09b (
    .a(al_6a408c69),
    .b(al_53bb123b[1]),
    .c(al_90a0fe97[0]),
    .o(al_18fbbb0f[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f13cf8f3 (
    .a(al_a4f25695),
    .b(al_1692563a[0]),
    .o(al_779bd70c[0]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_5f09fd11 (
    .a(al_cbeafa67[2]),
    .b(al_cbeafa67[4]),
    .c(al_cbeafa67[6]),
    .d(al_8932a489),
    .e(al_165f2734),
    .f(al_4c58e022),
    .o(al_b8b95ad1));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_76b61b55 (
    .a(al_b8b95ad1),
    .b(al_cbeafa67[0]),
    .c(al_90a0fe97[0]),
    .o(al_779bd70c[6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_23676f8a (
    .a(al_79090ab6),
    .b(al_41c9267e),
    .o(al_45d6e796[0]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_a96d8451 (
    .a(al_1ffff680),
    .o(al_56820b3e[2]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*B))"),
    .INIT(16'haa2a))
    al_8945ee1b (
    .a(al_2ccfdf18),
    .b(al_4ba8484b),
    .c(al_c5705f8a),
    .d(al_41c9267e),
    .o(al_56820b3e[6]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_546849bc (
    .a(al_79090ab6),
    .o(al_ff1cf72f));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_6f49a1ae (
    .a(al_be11f694),
    .b(al_ef9accde),
    .o(al_4ba8484b));
  AL_MAP_LUT3 #(
    .EQN("~(C*~B*A)"),
    .INIT(8'hdf))
    al_87850b48 (
    .a(al_be11f694),
    .b(al_ef9accde),
    .c(al_c58b049c),
    .o(al_f88e71cf));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    al_25583da2 (
    .a(al_f88e71cf),
    .b(al_4ba8484b),
    .o(al_a4f25695));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_942a42b7 (
    .a(al_a4f25695),
    .b(al_81cbac46[0]),
    .c(al_81c227e0[0]),
    .o(al_95504971[136]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_fa7e9066 (
    .a(al_2602b5cf[19]),
    .b(al_2602b5cf[29]),
    .c(al_2602b5cf[39]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_a2a57eb6));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_9d603b8f (
    .a(al_a4f25695),
    .b(al_a2a57eb6),
    .c(al_2602b5cf[9]),
    .d(al_81c227e0[0]),
    .o(al_95504971[64]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_7118a871 (
    .a(al_2602b5cf[18]),
    .b(al_2602b5cf[28]),
    .c(al_2602b5cf[38]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_9115a3ab));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_59795094 (
    .a(al_a4f25695),
    .b(al_9115a3ab),
    .c(al_2602b5cf[8]),
    .d(al_81c227e0[0]),
    .o(al_95504971[72]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_2579f1e0 (
    .a(al_2602b5cf[17]),
    .b(al_2602b5cf[27]),
    .c(al_2602b5cf[37]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_9b281de6));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_abb17067 (
    .a(al_a4f25695),
    .b(al_9b281de6),
    .c(al_2602b5cf[7]),
    .d(al_81c227e0[0]),
    .o(al_95504971[80]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_a9c00a5c (
    .a(al_2602b5cf[16]),
    .b(al_2602b5cf[26]),
    .c(al_2602b5cf[36]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_d3ca11f1));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_be61742f (
    .a(al_a4f25695),
    .b(al_d3ca11f1),
    .c(al_2602b5cf[6]),
    .d(al_81c227e0[0]),
    .o(al_95504971[88]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_4cc84fca (
    .a(al_2602b5cf[15]),
    .b(al_2602b5cf[25]),
    .c(al_2602b5cf[35]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_efe155a8));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_814281ed (
    .a(al_a4f25695),
    .b(al_efe155a8),
    .c(al_2602b5cf[5]),
    .d(al_81c227e0[0]),
    .o(al_95504971[96]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_5f4567b3 (
    .a(al_2602b5cf[14]),
    .b(al_2602b5cf[24]),
    .c(al_2602b5cf[34]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_f3fd3c4c));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_1d5e3651 (
    .a(al_a4f25695),
    .b(al_f3fd3c4c),
    .c(al_2602b5cf[4]),
    .d(al_81c227e0[0]),
    .o(al_95504971[104]));
  AL_MAP_LUT6 #(
    .EQN("(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*~(A)*~(D)+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*~(D)+~(((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E))*A*D+((F*C)*~(B)*~(E)+(F*C)*B*~(E)+~((F*C))*B*E+(F*C)*B*E)*A*D)"),
    .INIT(64'haaccaaf0aaccaa00))
    al_de45e384 (
    .a(al_2602b5cf[13]),
    .b(al_2602b5cf[23]),
    .c(al_2602b5cf[33]),
    .d(al_a26c7aae[1]),
    .e(al_a26c7aae[2]),
    .f(al_a26c7aae[3]),
    .o(al_8fe5c542));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_f305e2b9 (
    .a(al_a4f25695),
    .b(al_8fe5c542),
    .c(al_2602b5cf[3]),
    .d(al_81c227e0[0]),
    .o(al_95504971[112]));
  AL_DFF_0 al_5c31383c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_16ace516[27]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_dc65c0d1[21]));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_bfc3f610 (
    .a(1'b0),
    .o({al_dfdff5e7,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d30ddb3e (
    .a(al_e736aaf7[0]),
    .b(al_4f00db65),
    .c(al_dfdff5e7),
    .o({al_a45ee49d,al_9f02b6ff[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ae1798d1 (
    .a(al_e736aaf7[1]),
    .b(1'b0),
    .c(al_a45ee49d),
    .o({al_7de91657,al_9f02b6ff[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c75a04a5 (
    .a(al_e736aaf7[2]),
    .b(1'b0),
    .c(al_7de91657),
    .o({al_2fdead54,al_9f02b6ff[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_368a7200 (
    .a(al_e736aaf7[3]),
    .b(1'b0),
    .c(al_2fdead54),
    .o({al_73697ad3,al_9f02b6ff[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e587d1b7 (
    .a(al_e736aaf7[4]),
    .b(1'b0),
    .c(al_73697ad3),
    .o({al_482dfbbf,al_9f02b6ff[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_eda2fc21 (
    .a(al_e736aaf7[5]),
    .b(1'b0),
    .c(al_482dfbbf),
    .o({al_853f0be5,al_9f02b6ff[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e14a0894 (
    .a(al_e736aaf7[6]),
    .b(1'b0),
    .c(al_853f0be5),
    .o({al_b7fd68ad,al_9f02b6ff[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_13e1206 (
    .a(al_e736aaf7[7]),
    .b(1'b0),
    .c(al_b7fd68ad),
    .o({al_d323ca15,al_9f02b6ff[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c33ace2e (
    .a(al_e736aaf7[8]),
    .b(1'b0),
    .c(al_d323ca15),
    .o({al_7f632198,al_9f02b6ff[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_221d789 (
    .a(al_e736aaf7[9]),
    .b(1'b0),
    .c(al_7f632198),
    .o({al_35c78d09,al_9f02b6ff[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f4e51a40 (
    .a(al_e736aaf7[10]),
    .b(1'b0),
    .c(al_35c78d09),
    .o({al_6e02c90c,al_9f02b6ff[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2d80f51c (
    .a(al_e736aaf7[11]),
    .b(1'b0),
    .c(al_6e02c90c),
    .o({al_6f3fb610,al_9f02b6ff[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_381820ac (
    .a(al_e736aaf7[12]),
    .b(1'b0),
    .c(al_6f3fb610),
    .o({al_5f022649,al_9f02b6ff[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7f3d3266 (
    .a(al_e736aaf7[13]),
    .b(1'b0),
    .c(al_5f022649),
    .o({al_21c5d9e6,al_9f02b6ff[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9de7b955 (
    .a(al_e736aaf7[14]),
    .b(1'b0),
    .c(al_21c5d9e6),
    .o({al_312cedcc,al_9f02b6ff[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_12364d5a (
    .a(al_e736aaf7[15]),
    .b(1'b0),
    .c(al_312cedcc),
    .o({open_n3,al_9f02b6ff[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_c58b743a (
    .a(1'b0),
    .o({al_ba2fb587,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fc0cb8b9 (
    .a(al_a25915f6[0]),
    .b(1'b1),
    .c(al_ba2fb587),
    .o({al_f43a0c3c,al_b340bc6d[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c7aeaff9 (
    .a(al_a25915f6[1]),
    .b(1'b0),
    .c(al_f43a0c3c),
    .o({al_fd5b02e2,al_b340bc6d[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ac1c047a (
    .a(al_a25915f6[2]),
    .b(1'b0),
    .c(al_fd5b02e2),
    .o({al_9a41ae4f,al_b340bc6d[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d88c7f89 (
    .a(al_a25915f6[3]),
    .b(1'b0),
    .c(al_9a41ae4f),
    .o({al_b366bb58,al_b340bc6d[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8439005f (
    .a(al_a25915f6[4]),
    .b(1'b0),
    .c(al_b366bb58),
    .o({al_6784532f,al_b340bc6d[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7a819cc9 (
    .a(al_a25915f6[5]),
    .b(1'b0),
    .c(al_6784532f),
    .o({al_6c8827e1,al_b340bc6d[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_eda19a18 (
    .a(al_a25915f6[6]),
    .b(1'b0),
    .c(al_6c8827e1),
    .o({al_8a1c71af,al_b340bc6d[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e387b932 (
    .a(al_a25915f6[7]),
    .b(1'b0),
    .c(al_8a1c71af),
    .o({al_6d9415b,al_b340bc6d[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_92b1195c (
    .a(al_a25915f6[8]),
    .b(1'b0),
    .c(al_6d9415b),
    .o({al_e735abef,al_b340bc6d[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cd761d3 (
    .a(al_a25915f6[9]),
    .b(1'b0),
    .c(al_e735abef),
    .o({al_2a364bea,al_b340bc6d[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_680a1630 (
    .a(al_a25915f6[10]),
    .b(1'b0),
    .c(al_2a364bea),
    .o({al_1cc7635e,al_b340bc6d[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f3673a14 (
    .a(al_a25915f6[11]),
    .b(1'b0),
    .c(al_1cc7635e),
    .o({al_c4e50727,al_b340bc6d[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_72da9815 (
    .a(al_a25915f6[12]),
    .b(1'b0),
    .c(al_c4e50727),
    .o({al_aa8528c4,al_b340bc6d[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1ec9b5f3 (
    .a(al_a25915f6[13]),
    .b(1'b0),
    .c(al_aa8528c4),
    .o({al_12af440,al_b340bc6d[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_25d1b1bd (
    .a(al_a25915f6[14]),
    .b(1'b0),
    .c(al_12af440),
    .o({al_174c5495,al_b340bc6d[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_be00d667 (
    .a(al_a25915f6[15]),
    .b(1'b0),
    .c(al_174c5495),
    .o({open_n7,al_b340bc6d[15]}));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~A*~(E*D*C)))"),
    .INIT(32'h32222222))
    al_312d3037 (
    .a(al_45d2984c),
    .b(al_eec1ba11),
    .c(al_9ffa2c81[0]),
    .d(al_9ffa2c81[1]),
    .e(al_9ffa2c81[2]),
    .o(al_855245d9));
  AL_DFF_0 al_73efcb1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_855245d9),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_45d2984c));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(C*B)))"),
    .INIT(16'h00d5))
    al_72c42292 (
    .a(al_9120ce24),
    .b(al_81cbac46[0]),
    .c(al_81c227e0[0]),
    .d(al_eec1ba11),
    .o(al_5a67a09b[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_10b02ae1 (
    .a(al_eec1ba11),
    .b(al_9ffa2c81[0]),
    .o(al_5a67a09b[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_de147a6f (
    .a(al_eec1ba11),
    .b(al_9ffa2c81[1]),
    .o(al_5a67a09b[2]));
  AL_MAP_LUT6 #(
    .EQN("~(~(~F*E*D*~C)*~(B*~A))"),
    .INIT(64'h444444444f444444))
    al_20d98997 (
    .a(al_147f1ed5[0]),
    .b(al_147f1ed5[1]),
    .c(al_2e186afc[0]),
    .d(al_2e186afc[1]),
    .e(al_2e186afc[2]),
    .f(al_2e186afc[3]),
    .o(al_ac2c2542[0]));
  AL_MAP_LUT6 #(
    .EQN("~(~(~F*E*D*~C)*~(B*A))"),
    .INIT(64'h888888888f888888))
    al_c5fd94dc (
    .a(al_147f1ed5[0]),
    .b(al_147f1ed5[1]),
    .c(al_2e186afc[0]),
    .d(al_2e186afc[1]),
    .e(al_2e186afc[2]),
    .f(al_2e186afc[3]),
    .o(al_ac2c2542[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_976f546e (
    .a(al_147f1ed5[0]),
    .b(al_147f1ed5[1]),
    .o(al_68e325c6));
  AL_MAP_LUT5 #(
    .EQN("~((D*C*A)*~(E)*~(B)+(D*C*A)*E*~(B)+~((D*C*A))*E*B+(D*C*A)*E*B)"),
    .INIT(32'h1333dfff))
    al_475eaa37 (
    .a(al_58bba036),
    .b(al_2e186afc[0]),
    .c(al_1d853c9a[0]),
    .d(al_1d853c9a[1]),
    .e(al_898823b1),
    .o(al_66c80cd2));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hcccc000fff00aaaa))
    al_c867cb (
    .a(al_66c80cd2),
    .b(al_e4885785),
    .c(al_58ef9f1a),
    .d(al_2e186afc[0]),
    .e(al_2e186afc[1]),
    .f(al_2e186afc[2]),
    .o(al_7f9da669));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_cddc0810 (
    .a(al_7f9da669),
    .b(al_2e186afc[3]),
    .o(al_c3b79934[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_cff20409 (
    .a(al_147f1ed5[0]),
    .b(al_147f1ed5[1]),
    .c(al_2e186afc[0]),
    .o(al_e4885785));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_af07efb3 (
    .a(al_1d853c9a[2]),
    .b(al_1d853c9a[3]),
    .o(al_1495678c));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_17b52864 (
    .a(al_1495678c),
    .b(al_1d853c9a[0]),
    .c(al_1d853c9a[1]),
    .o(al_a6bf875b));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfdc1))
    al_d33ac7c0 (
    .a(al_a6bf875b),
    .b(al_2e186afc[0]),
    .c(al_2e186afc[1]),
    .d(al_898823b1),
    .o(al_a807e4d3));
  AL_MAP_LUT5 #(
    .EQN("(~E*(~A*~((C*~B))*~(D)+~A*(C*~B)*~(D)+~(~A)*(C*~B)*D+~A*(C*~B)*D))"),
    .INIT(32'h00003055))
    al_7bdbbef0 (
    .a(al_a807e4d3),
    .b(al_e4885785),
    .c(al_2e186afc[1]),
    .d(al_2e186afc[2]),
    .e(al_2e186afc[3]),
    .o(al_c3b79934[1]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E))"),
    .INIT(64'h0000000033fff00a))
    al_bab5e150 (
    .a(al_a6bf875b),
    .b(al_e4885785),
    .c(al_2e186afc[0]),
    .d(al_2e186afc[1]),
    .e(al_2e186afc[2]),
    .f(al_2e186afc[3]),
    .o(al_c3b79934[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_907c1c68 (
    .a(al_e4885785),
    .b(al_2e186afc[1]),
    .c(al_2e186afc[2]),
    .d(al_2e186afc[3]),
    .o(al_c3b79934[3]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*~B*~A)"),
    .INIT(64'h1000000000000000))
    al_7fb4c7e7 (
    .a(al_eec1ba11),
    .b(al_a25915f6[0]),
    .c(al_a25915f6[1]),
    .d(al_a25915f6[2]),
    .e(al_a25915f6[3]),
    .f(al_a25915f6[4]),
    .o(al_713543ac));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_772adeab (
    .a(al_a25915f6[5]),
    .b(al_a25915f6[6]),
    .c(al_a25915f6[7]),
    .d(al_a25915f6[8]),
    .o(al_c0d8b545));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_a1f77943 (
    .a(al_c0d8b545),
    .b(al_a25915f6[9]),
    .c(al_a25915f6[10]),
    .d(al_a25915f6[11]),
    .e(al_a25915f6[12]),
    .o(al_24009166));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_c643bf9b (
    .a(al_24009166),
    .b(al_713543ac),
    .c(al_a25915f6[13]),
    .d(al_a25915f6[14]),
    .e(al_a25915f6[15]),
    .o(al_ca978bef));
  AL_DFF_0 al_f5aa8655 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ca978bef),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f00db65));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*B)*~(~E*~D*A))"),
    .INIT(32'hc0c0c0ea))
    al_88fb293d (
    .a(al_58bba036),
    .b(al_6d33eaeb),
    .c(al_20ae9484),
    .d(al_1d853c9a[0]),
    .e(al_1d853c9a[1]),
    .o(al_dc674b57));
  AL_DFF_0 al_8b8928f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dc674b57),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eec1ba11));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_498e89bf (
    .a(al_e736aaf7[0]),
    .b(al_e736aaf7[1]),
    .c(al_e736aaf7[2]),
    .d(al_e736aaf7[3]),
    .o(al_a3c61604));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_82ecc310 (
    .a(al_e736aaf7[8]),
    .b(al_e736aaf7[9]),
    .c(al_e736aaf7[10]),
    .d(al_e736aaf7[11]),
    .o(al_7fdd8f7a));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_578b13be (
    .a(al_7fdd8f7a),
    .b(al_e736aaf7[12]),
    .c(al_e736aaf7[13]),
    .d(al_e736aaf7[14]),
    .e(al_e736aaf7[15]),
    .o(al_b16882ef));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_c410bc44 (
    .a(al_b16882ef),
    .b(al_a3c61604),
    .c(al_e736aaf7[4]),
    .d(al_e736aaf7[5]),
    .e(al_e736aaf7[6]),
    .f(al_e736aaf7[7]),
    .o(al_fa46dbba));
  AL_DFF_0 al_bd024de2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fa46dbba),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d33eaeb));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_d0bdb7fe (
    .a(al_a25915f6[4]),
    .b(al_a25915f6[5]),
    .c(al_a25915f6[6]),
    .d(al_a25915f6[7]),
    .o(al_370abec1));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_305a8ea3 (
    .a(al_370abec1),
    .b(al_a25915f6[0]),
    .c(al_a25915f6[1]),
    .d(al_a25915f6[2]),
    .e(al_a25915f6[3]),
    .o(al_15b509ab));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_9e57fb23 (
    .a(al_a25915f6[8]),
    .b(al_a25915f6[9]),
    .c(al_a25915f6[10]),
    .d(al_a25915f6[11]),
    .o(al_6255d7f7));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_de85d75d (
    .a(al_15b509ab),
    .b(al_6255d7f7),
    .c(al_a25915f6[12]),
    .d(al_a25915f6[13]),
    .e(al_a25915f6[14]),
    .f(al_a25915f6[15]),
    .o(al_3f6a9f97));
  AL_DFF_0 al_78eb51c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3f6a9f97),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_20ae9484));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_ada188f5 (
    .a(al_b5a5e144),
    .b(al_eec1ba11),
    .o(al_1fe9b96a));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_2b9dbaee (
    .a(al_2e186afc[0]),
    .b(al_2e186afc[1]),
    .c(al_2e186afc[2]),
    .d(al_2e186afc[3]),
    .o(al_afe8a6f9));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_1a222607 (
    .a(al_2e186afc[0]),
    .b(al_2e186afc[1]),
    .c(al_898823b1),
    .o(al_18aca87e));
  AL_MAP_LUT5 #(
    .EQN("~(~B*(A*~(C)*D*~(E)+~(A)*C*~(D)*E+A*C*~(D)*E+A*~(C)*D*E))"),
    .INIT(32'hfdcffdff))
    al_c503097e (
    .a(al_58ef9f1a),
    .b(al_2e186afc[0]),
    .c(al_2e186afc[1]),
    .d(al_2e186afc[2]),
    .e(al_898823b1),
    .o(al_f57af6b4));
  AL_MAP_LUT5 #(
    .EQN("(A*C*~((~D*B))*~(E)+A*~(C)*(~D*B)*~(E)+A*C*(~D*B)*~(E)+~(A)*C*~((~D*B))*E+A*C*~((~D*B))*E+~(A)*C*(~D*B)*E+A*C*(~D*B)*E)"),
    .INIT(32'hf0f0a0a8))
    al_ca0329c5 (
    .a(al_f57af6b4),
    .b(al_18aca87e),
    .c(al_a082bc48),
    .d(al_2e186afc[2]),
    .e(al_2e186afc[3]),
    .o(al_154c9279));
  AL_DFF_0 al_896fac55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_154c9279),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a082bc48));
  AL_DFF_0 al_94f5bdb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_68e325c6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58b049c));
  AL_DFF_0 al_a5cc64a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_afe8a6f9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b38e0f3));
  AL_DFF_0 al_1a9d5482 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(init_calib_complete),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b2bde781));
  AL_MAP_LUT6 #(
    .EQN("(~E*A*(D*~((C*B))*~(F)+D*(C*B)*~(F)+~(D)*(C*B)*F+D*(C*B)*F))"),
    .INIT(64'h000080800000aa00))
    al_f8b70cd3 (
    .a(al_58bba036),
    .b(al_6d33eaeb),
    .c(al_20ae9484),
    .d(al_b2bde781),
    .e(al_1d853c9a[0]),
    .f(al_1d853c9a[1]),
    .o(al_fc9b7dfa));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(~D*C*A))"),
    .INIT(16'hccec))
    al_ae0a4670 (
    .a(al_7959b11f),
    .b(al_fc9b7dfa),
    .c(al_1495678c),
    .d(al_1d853c9a[0]),
    .o(al_da91be3[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_20e04693 (
    .a(al_1d853c9a[2]),
    .b(al_1d853c9a[3]),
    .o(al_58bba036));
  AL_MAP_LUT5 #(
    .EQN("~(A*~(C*(~(B)*D*~(E)+B*D*~(E)+~(B)*~(D)*E)))"),
    .INIT(32'h5575f555))
    al_efdb0add (
    .a(al_484f859d),
    .b(al_22ec870),
    .c(al_58bba036),
    .d(al_1d853c9a[0]),
    .e(al_1d853c9a[1]),
    .o(al_da91be3[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_5f73c200 (
    .a(al_2e186afc[0]),
    .b(al_2e186afc[1]),
    .o(al_90876008));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_676bcf73 (
    .a(al_90876008),
    .b(al_2e186afc[2]),
    .c(al_2e186afc[3]),
    .o(al_7959b11f));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    al_a8e10be1 (
    .a(al_45d2984c),
    .b(al_6d33eaeb),
    .c(al_20ae9484),
    .d(al_69c9761a),
    .o(al_22ec870));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfffffff3f005ffff))
    al_6085d733 (
    .a(al_7959b11f),
    .b(al_b2bde781),
    .c(al_1d853c9a[0]),
    .d(al_1d853c9a[1]),
    .e(al_1d853c9a[2]),
    .f(al_1d853c9a[3]),
    .o(al_484f859d));
  AL_MAP_LUT6 #(
    .EQN("(~((C*B*A))*~(D)*~(E)*~(F)+(C*B*A)*~(D)*~(E)*~(F)+~((C*B*A))*D*~(E)*~(F)+(C*B*A)*D*~(E)*~(F)+~((C*B*A))*~(D)*E*~(F)+~((C*B*A))*D*E*F+(C*B*A)*D*E*F)"),
    .INIT(64'hff000000007fffff))
    al_3c1d9ac9 (
    .a(al_6d33eaeb),
    .b(al_20ae9484),
    .c(al_69c9761a),
    .d(al_1d853c9a[0]),
    .e(al_1d853c9a[1]),
    .f(al_1d853c9a[2]),
    .o(al_9b835e77));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_f713f93b (
    .a(al_9b835e77),
    .b(al_1d853c9a[3]),
    .o(al_da91be3[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_6cc968c8 (
    .a(al_1495678c),
    .b(al_1d853c9a[0]),
    .c(al_1d853c9a[1]),
    .o(al_da91be3[3]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~(A*~(C*B))))"),
    .INIT(32'h00ff002a))
    al_5a357efd (
    .a(al_9120ce24),
    .b(al_81cbac46[0]),
    .c(al_81c227e0[0]),
    .d(al_eec1ba11),
    .e(al_69c9761a),
    .o(al_67ffb718));
  AL_DFF_0 al_5bee8c8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_67ffb718),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_69c9761a));
  AL_DFF_0 al_3c9ddd59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a67a09b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9ffa2c81[0]));
  AL_DFF_0 al_63972aa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a67a09b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9ffa2c81[1]));
  AL_DFF_0 al_891ca9ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a67a09b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9ffa2c81[2]));
  AL_DFF_0 al_58b38b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ac2c2542[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_147f1ed5[0]));
  AL_DFF_0 al_7bf7a94f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ac2c2542[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_147f1ed5[1]));
  AL_DFF_0 al_419dcfef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3b79934[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_2e186afc[0]));
  AL_DFF_0 al_53dac869 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3b79934[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_2e186afc[1]));
  AL_DFF_0 al_e9bc83fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3b79934[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_2e186afc[2]));
  AL_DFF_0 al_48c2373e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3b79934[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_2e186afc[3]));
  AL_DFF_0 al_aa10050d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[0]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[0]));
  AL_DFF_0 al_e95c0ca0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[1]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[1]));
  AL_DFF_0 al_dbbb0d1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[2]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[2]));
  AL_DFF_0 al_2915007b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[3]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[3]));
  AL_DFF_0 al_41e6b71d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[4]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[4]));
  AL_DFF_0 al_e72a7d2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[5]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[5]));
  AL_DFF_0 al_17db8492 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[6]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[6]));
  AL_DFF_0 al_c6cfe970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[7]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[7]));
  AL_DFF_0 al_238b8cf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[8]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[8]));
  AL_DFF_0 al_99d2dec7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[9]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[9]));
  AL_DFF_0 al_e75aa1b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[10]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[10]));
  AL_DFF_0 al_91bd4b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[11]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[11]));
  AL_DFF_0 al_772ab2db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[12]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[12]));
  AL_DFF_0 al_e660c741 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[13]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[13]));
  AL_DFF_0 al_3bb9985 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[14]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[14]));
  AL_DFF_0 al_38ddb4e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f02b6ff[15]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_e736aaf7[15]));
  AL_DFF_0 al_b5acc303 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[0]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[0]));
  AL_DFF_0 al_5aaf5e11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[1]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[1]));
  AL_DFF_0 al_afd69be8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[2]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[2]));
  AL_DFF_0 al_307ad82e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[3]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[3]));
  AL_DFF_0 al_dd63798f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[4]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[4]));
  AL_DFF_0 al_802a0462 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[5]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[5]));
  AL_DFF_0 al_40d7e92e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[6]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[6]));
  AL_DFF_0 al_90fb9563 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[7]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[7]));
  AL_DFF_0 al_7f2545ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[8]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[8]));
  AL_DFF_0 al_5987faf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[9]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[9]));
  AL_DFF_0 al_dcc3f9d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[10]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[10]));
  AL_DFF_0 al_6a2beee7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[11]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[11]));
  AL_DFF_0 al_4f579e45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[12]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[12]));
  AL_DFF_0 al_c44e07e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[13]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[13]));
  AL_DFF_0 al_5eecf3eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[14]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[14]));
  AL_DFF_0 al_907dab73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b340bc6d[15]),
    .en(1'b1),
    .sr(~al_1fe9b96a),
    .ss(1'b0),
    .q(al_a25915f6[15]));
  AL_DFF_0 al_b0dad259 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_da91be3[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_1d853c9a[0]));
  AL_DFF_0 al_944314b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_da91be3[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_1d853c9a[1]));
  AL_DFF_0 al_f17b1378 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_da91be3[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_1d853c9a[2]));
  AL_DFF_0 al_b2ba202e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_da91be3[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_1d853c9a[3]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*~B*~A)"),
    .INIT(16'hfffe))
    al_d4c6287d (
    .a(al_8d73b4c8[0]),
    .b(al_8d73b4c8[1]),
    .c(al_8d73b4c8[2]),
    .d(al_8d73b4c8[3]),
    .o(al_432340bb));
  AL_DFF_0 al_c4f3a242 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_432340bb),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5bb559f0));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*~B*~A)"),
    .INIT(16'hfffe))
    al_667ca070 (
    .a(al_f4295ad6[0]),
    .b(al_f4295ad6[1]),
    .c(al_f4295ad6[2]),
    .d(al_f4295ad6[3]),
    .o(al_ee2d8b77));
  AL_DFF_0 al_f6d50335 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ee2d8b77),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_3f592f2c));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    al_152dda11 (
    .a(al_887856fc[0]),
    .b(al_5bb559f0),
    .c(al_3f592f2c),
    .o(al_a8d985cf[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    al_85b42c77 (
    .a(al_b4c6b3bd),
    .b(al_d50c8b50),
    .c(al_5bb559f0),
    .d(al_3f592f2c),
    .o(al_a8d985cf[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    al_6de7a837 (
    .a(al_ef78cbcb),
    .b(al_a70d3eb4),
    .c(al_5bb559f0),
    .d(al_3f592f2c),
    .o(al_a8d985cf[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    al_cb19be33 (
    .a(al_887856fc[3]),
    .b(al_5bb559f0),
    .c(al_3f592f2c),
    .o(al_a8d985cf[3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(~D*B)))"),
    .INIT(16'ha028))
    al_e0f0942 (
    .a(al_d99aae4d[0]),
    .b(al_5e053069[0]),
    .c(al_5e053069[1]),
    .d(al_f4295ad6[0]),
    .o(al_6c3719db[1]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_1bf768bf (
    .a(al_55232c98),
    .b(al_d99aae4d[0]),
    .c(al_5e053069[2]),
    .d(al_5e053069[3]),
    .e(al_5e053069[4]),
    .o(al_6c3719db[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_e0e83ae9 (
    .a(al_524ab3e2),
    .b(al_d99aae4d[0]),
    .c(al_5e053069[5]),
    .d(al_5e053069[6]),
    .e(al_5e053069[7]),
    .o(al_6c3719db[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(~D*B)))"),
    .INIT(16'ha028))
    al_5f6248df (
    .a(al_d99aae4d[1]),
    .b(al_d07272c1[0]),
    .c(al_d07272c1[1]),
    .d(al_f4295ad6[1]),
    .o(al_fd291354[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_3fa78416 (
    .a(al_be5b15b0),
    .b(al_d99aae4d[1]),
    .c(al_d07272c1[4]),
    .o(al_fd291354[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_b5be0109 (
    .a(al_685b247),
    .b(al_d99aae4d[1]),
    .c(al_d07272c1[5]),
    .d(al_d07272c1[6]),
    .e(al_d07272c1[7]),
    .o(al_fd291354[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(~D*B)))"),
    .INIT(16'ha028))
    al_7d1c7af5 (
    .a(al_d99aae4d[2]),
    .b(al_582cdf5[0]),
    .c(al_582cdf5[1]),
    .d(al_f4295ad6[2]),
    .o(al_7861e435[1]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_a7ea0cbe (
    .a(al_698dfed0),
    .b(al_d99aae4d[2]),
    .c(al_582cdf5[2]),
    .d(al_582cdf5[3]),
    .e(al_582cdf5[4]),
    .o(al_7861e435[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_e1d77fff (
    .a(al_1223a962),
    .b(al_d99aae4d[2]),
    .c(al_582cdf5[5]),
    .d(al_582cdf5[6]),
    .e(al_582cdf5[7]),
    .o(al_7861e435[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(~D*B)))"),
    .INIT(16'ha028))
    al_1ae5d1c5 (
    .a(al_d99aae4d[3]),
    .b(al_a3070745[0]),
    .c(al_a3070745[1]),
    .d(al_f4295ad6[3]),
    .o(al_9c26f92c[1]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_f9f3027e (
    .a(al_2d260a04),
    .b(al_d99aae4d[3]),
    .c(al_a3070745[2]),
    .d(al_a3070745[3]),
    .e(al_a3070745[4]),
    .o(al_9c26f92c[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_8ad5a94d (
    .a(al_12563419),
    .b(al_d99aae4d[3]),
    .c(al_a3070745[5]),
    .d(al_a3070745[6]),
    .e(al_a3070745[7]),
    .o(al_9c26f92c[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_8b332183 (
    .a(al_d99aae4d[0]),
    .b(al_5e053069[0]),
    .c(al_f4295ad6[0]),
    .o(al_6c3719db[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_5cad7bc3 (
    .a(al_a76392f),
    .b(al_6c3719db[5]),
    .c(al_6c3719db[6]),
    .d(al_6c3719db[8]),
    .o(al_82fe8ddf[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_aab16c4f (
    .a(al_5e053069[0]),
    .b(al_5e053069[1]),
    .c(al_f4295ad6[0]),
    .o(al_55232c98));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_7025c93d (
    .a(al_55232c98),
    .b(al_d99aae4d[0]),
    .c(al_5e053069[2]),
    .o(al_6c3719db[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_d85ad5c9 (
    .a(al_55232c98),
    .b(al_d99aae4d[0]),
    .c(al_5e053069[2]),
    .d(al_5e053069[3]),
    .o(al_6c3719db[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_a6f106a7 (
    .a(al_55232c98),
    .b(al_5e053069[2]),
    .c(al_5e053069[3]),
    .d(al_5e053069[4]),
    .o(al_524ab3e2));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_380cb216 (
    .a(al_524ab3e2),
    .b(al_d99aae4d[0]),
    .c(al_5e053069[5]),
    .o(al_6c3719db[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_3377c138 (
    .a(al_524ab3e2),
    .b(al_d99aae4d[0]),
    .c(al_5e053069[5]),
    .d(al_5e053069[6]),
    .o(al_6c3719db[6]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_f558096c (
    .a(al_524ab3e2),
    .b(al_d99aae4d[0]),
    .c(al_5e053069[5]),
    .d(al_5e053069[6]),
    .e(al_5e053069[7]),
    .f(al_5e053069[8]),
    .o(al_6c3719db[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_ca45a0af (
    .a(al_6c3719db[2]),
    .b(al_6c3719db[3]),
    .c(al_6c3719db[0]),
    .d(al_5e053069[1]),
    .e(al_5e053069[4]),
    .f(al_5e053069[7]),
    .o(al_a76392f));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_8d9893f8 (
    .a(al_d99aae4d[1]),
    .b(al_d07272c1[0]),
    .c(al_f4295ad6[1]),
    .o(al_fd291354[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_59988485 (
    .a(al_fd291354[5]),
    .b(al_fd291354[6]),
    .c(al_fd291354[8]),
    .d(al_5ece979a),
    .o(al_82fe8ddf[1]));
  AL_MAP_LUT5 #(
    .EQN("(A*(D@(~E*C*B)))"),
    .INIT(32'haa002a80))
    al_a9ff11df (
    .a(al_d99aae4d[1]),
    .b(al_d07272c1[0]),
    .c(al_d07272c1[1]),
    .d(al_d07272c1[2]),
    .e(al_f4295ad6[1]),
    .o(al_fd291354[2]));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    al_b4ac08e1 (
    .a(al_d07272c1[0]),
    .b(al_d07272c1[1]),
    .c(al_d07272c1[2]),
    .d(al_d07272c1[3]),
    .e(al_f4295ad6[1]),
    .o(al_be5b15b0));
  AL_MAP_LUT6 #(
    .EQN("(A*(E@(~F*D*C*B)))"),
    .INIT(64'haaaa00002aaa8000))
    al_eb241298 (
    .a(al_d99aae4d[1]),
    .b(al_d07272c1[0]),
    .c(al_d07272c1[1]),
    .d(al_d07272c1[2]),
    .e(al_d07272c1[3]),
    .f(al_f4295ad6[1]),
    .o(al_fd291354[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_c5a612e4 (
    .a(al_be5b15b0),
    .b(al_d07272c1[4]),
    .o(al_685b247));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_7460c3c3 (
    .a(al_685b247),
    .b(al_d99aae4d[1]),
    .c(al_d07272c1[5]),
    .o(al_fd291354[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_bfe40d51 (
    .a(al_685b247),
    .b(al_d99aae4d[1]),
    .c(al_d07272c1[5]),
    .d(al_d07272c1[6]),
    .o(al_fd291354[6]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_fde471f8 (
    .a(al_685b247),
    .b(al_d99aae4d[1]),
    .c(al_d07272c1[5]),
    .d(al_d07272c1[6]),
    .e(al_d07272c1[7]),
    .f(al_d07272c1[8]),
    .o(al_fd291354[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_fa062b04 (
    .a(al_fd291354[3]),
    .b(al_fd291354[2]),
    .c(al_fd291354[0]),
    .d(al_d07272c1[1]),
    .e(al_d07272c1[4]),
    .f(al_d07272c1[7]),
    .o(al_5ece979a));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_e905d6a8 (
    .a(al_d99aae4d[2]),
    .b(al_582cdf5[0]),
    .c(al_f4295ad6[2]),
    .o(al_7861e435[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_ef4b9563 (
    .a(al_e29cf77),
    .b(al_7861e435[5]),
    .c(al_7861e435[6]),
    .d(al_7861e435[8]),
    .o(al_82fe8ddf[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_f76be24c (
    .a(al_582cdf5[0]),
    .b(al_582cdf5[1]),
    .c(al_f4295ad6[2]),
    .o(al_698dfed0));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_11c6305c (
    .a(al_698dfed0),
    .b(al_d99aae4d[2]),
    .c(al_582cdf5[2]),
    .o(al_7861e435[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_55786179 (
    .a(al_698dfed0),
    .b(al_d99aae4d[2]),
    .c(al_582cdf5[2]),
    .d(al_582cdf5[3]),
    .o(al_7861e435[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_c98141c1 (
    .a(al_698dfed0),
    .b(al_582cdf5[2]),
    .c(al_582cdf5[3]),
    .d(al_582cdf5[4]),
    .o(al_1223a962));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_4bcd3c1 (
    .a(al_1223a962),
    .b(al_d99aae4d[2]),
    .c(al_582cdf5[5]),
    .o(al_7861e435[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_e53f2b8d (
    .a(al_1223a962),
    .b(al_d99aae4d[2]),
    .c(al_582cdf5[5]),
    .d(al_582cdf5[6]),
    .o(al_7861e435[6]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_49567385 (
    .a(al_1223a962),
    .b(al_d99aae4d[2]),
    .c(al_582cdf5[5]),
    .d(al_582cdf5[6]),
    .e(al_582cdf5[7]),
    .f(al_582cdf5[8]),
    .o(al_7861e435[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_fbc38ae4 (
    .a(al_7861e435[2]),
    .b(al_7861e435[3]),
    .c(al_7861e435[0]),
    .d(al_582cdf5[1]),
    .e(al_582cdf5[4]),
    .f(al_582cdf5[7]),
    .o(al_e29cf77));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_43d74899 (
    .a(al_d99aae4d[3]),
    .b(al_a3070745[0]),
    .c(al_f4295ad6[3]),
    .o(al_9c26f92c[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_248e7fa4 (
    .a(al_bc808160),
    .b(al_9c26f92c[5]),
    .c(al_9c26f92c[6]),
    .d(al_9c26f92c[8]),
    .o(al_82fe8ddf[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_ceb1725f (
    .a(al_a3070745[0]),
    .b(al_a3070745[1]),
    .c(al_f4295ad6[3]),
    .o(al_2d260a04));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_428affd2 (
    .a(al_2d260a04),
    .b(al_d99aae4d[3]),
    .c(al_a3070745[2]),
    .o(al_9c26f92c[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_38efa311 (
    .a(al_2d260a04),
    .b(al_d99aae4d[3]),
    .c(al_a3070745[2]),
    .d(al_a3070745[3]),
    .o(al_9c26f92c[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_6f35063d (
    .a(al_2d260a04),
    .b(al_a3070745[2]),
    .c(al_a3070745[3]),
    .d(al_a3070745[4]),
    .o(al_12563419));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_84bb8c9 (
    .a(al_12563419),
    .b(al_d99aae4d[3]),
    .c(al_a3070745[5]),
    .o(al_9c26f92c[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_403a3993 (
    .a(al_12563419),
    .b(al_d99aae4d[3]),
    .c(al_a3070745[5]),
    .d(al_a3070745[6]),
    .o(al_9c26f92c[6]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_5e04b5e6 (
    .a(al_12563419),
    .b(al_d99aae4d[3]),
    .c(al_a3070745[5]),
    .d(al_a3070745[6]),
    .e(al_a3070745[7]),
    .f(al_a3070745[8]),
    .o(al_9c26f92c[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_4b0ab362 (
    .a(al_9c26f92c[2]),
    .b(al_9c26f92c[3]),
    .c(al_9c26f92c[0]),
    .d(al_a3070745[1]),
    .e(al_a3070745[4]),
    .f(al_a3070745[7]),
    .o(al_bc808160));
  AL_DFF_0 al_340b0431 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a8d985cf[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d99aae4d[0]));
  AL_DFF_0 al_bafd617b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a8d985cf[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d99aae4d[1]));
  AL_DFF_0 al_20ab8ef3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a8d985cf[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d99aae4d[2]));
  AL_DFF_0 al_fdbabb6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a8d985cf[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d99aae4d[3]));
  AL_DFF_0 al_31e8146a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[0]));
  AL_DFF_0 al_ac4f33ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[1]));
  AL_DFF_0 al_741ed5e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[2]));
  AL_DFF_0 al_9cbbaf45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[3]));
  AL_DFF_0 al_6e8eb6f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[4]));
  AL_DFF_0 al_b796a9d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[5]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[5]));
  AL_DFF_0 al_6ad893fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[6]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[6]));
  AL_DFF_0 al_a4c66444 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[7]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[7]));
  AL_DFF_0 al_c3513eba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c3719db[8]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_5e053069[8]));
  AL_DFF_0 al_4371e38e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[0]));
  AL_DFF_0 al_512606a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[1]));
  AL_DFF_0 al_11e22bfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[2]));
  AL_DFF_0 al_2f88fd22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[3]));
  AL_DFF_0 al_611c418b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[4]));
  AL_DFF_0 al_c45af13b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[5]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[5]));
  AL_DFF_0 al_bd4fb3cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[6]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[6]));
  AL_DFF_0 al_8f845d3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[7]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[7]));
  AL_DFF_0 al_6a8d53a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd291354[8]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d07272c1[8]));
  AL_DFF_0 al_1cd64a6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[0]));
  AL_DFF_0 al_c4cdfa6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[1]));
  AL_DFF_0 al_13e5ea1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[2]));
  AL_DFF_0 al_210f3e5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[3]));
  AL_DFF_0 al_2ef8d379 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[4]));
  AL_DFF_0 al_4a5cf4cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[5]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[5]));
  AL_DFF_0 al_dc1c4e7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[6]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[6]));
  AL_DFF_0 al_f67a459d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[7]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[7]));
  AL_DFF_0 al_f86b4123 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7861e435[8]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_582cdf5[8]));
  AL_DFF_0 al_615a7772 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[0]));
  AL_DFF_0 al_3c119cd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[1]));
  AL_DFF_0 al_1d6689fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[2]));
  AL_DFF_0 al_cb5cb9eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[3]));
  AL_DFF_0 al_40c587fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[4]));
  AL_DFF_0 al_847367e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[5]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[5]));
  AL_DFF_0 al_32d3b212 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[6]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[6]));
  AL_DFF_0 al_9b7507d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[7]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[7]));
  AL_DFF_0 al_d2b35e8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c26f92c[8]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_a3070745[8]));
  AL_DFF_0 al_20157043 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_82fe8ddf[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_f4295ad6[0]));
  AL_DFF_0 al_f240c697 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_82fe8ddf[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_f4295ad6[1]));
  AL_DFF_0 al_7a8994b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_82fe8ddf[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_f4295ad6[2]));
  AL_DFF_0 al_93167cab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_82fe8ddf[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_f4295ad6[3]));
  AL_DFF_0 al_99628b74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_93b093ad[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_92b55720[0]));
  AL_DFF_0 al_e87b27d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_93b093ad[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_92b55720[1]));
  AL_DFF_0 al_59580697 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_93b093ad[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_92b55720[2]));
  AL_DFF_0 al_913895db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_93b093ad[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_92b55720[3]));
  AL_DFF_0 al_bf8ad937 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[0]));
  AL_DFF_0 al_489f71a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[1]));
  AL_DFF_0 al_a979823b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[2]));
  AL_DFF_0 al_1f4b7198 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[3]));
  AL_DFF_0 al_1165a3d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[4]));
  AL_DFF_0 al_14b23f7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[5]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[5]));
  AL_DFF_0 al_4368f40c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[6]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[6]));
  AL_DFF_0 al_4c9d6ae4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[7]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[7]));
  AL_DFF_0 al_47702388 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dedaebcb[8]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_52b895b5[8]));
  AL_DFF_0 al_1a02b69d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[0]));
  AL_DFF_0 al_5ac46c1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[1]));
  AL_DFF_0 al_b8a5931e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[2]));
  AL_DFF_0 al_e114f199 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[3]));
  AL_DFF_0 al_2d4d011e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[4]));
  AL_DFF_0 al_b169d767 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[5]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[5]));
  AL_DFF_0 al_c175092e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[6]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[6]));
  AL_DFF_0 al_51a829e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[7]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[7]));
  AL_DFF_0 al_6d259079 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6fe26a79[8]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_bd6aead3[8]));
  AL_DFF_0 al_55e754da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[0]));
  AL_DFF_0 al_19514e03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[1]));
  AL_DFF_0 al_9b59f31b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[2]));
  AL_DFF_0 al_7b763d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[3]));
  AL_DFF_0 al_428b9c74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[4]));
  AL_DFF_0 al_95f52619 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[5]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[5]));
  AL_DFF_0 al_11b4a316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[6]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[6]));
  AL_DFF_0 al_e14585c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[7]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[7]));
  AL_DFF_0 al_8d35080b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_910cb5e3[8]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_febad4d6[8]));
  AL_DFF_0 al_6ae4c92a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[0]));
  AL_DFF_0 al_e77d9788 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[1]));
  AL_DFF_0 al_ba01b795 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[2]));
  AL_DFF_0 al_b3179e06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[3]));
  AL_DFF_0 al_1df8d69b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[4]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[4]));
  AL_DFF_0 al_4a71acce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[5]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[5]));
  AL_DFF_0 al_359739f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[6]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[6]));
  AL_DFF_0 al_549e8bef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[7]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[7]));
  AL_DFF_0 al_3e492e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b9547a0[8]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c57192d3[8]));
  AL_DFF_0 al_a3a93eae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e39e8b51[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_8d73b4c8[0]));
  AL_DFF_0 al_d596e90a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e39e8b51[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_8d73b4c8[1]));
  AL_DFF_0 al_ab6b74ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e39e8b51[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_8d73b4c8[2]));
  AL_DFF_0 al_a0cb4aa3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e39e8b51[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_8d73b4c8[3]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_498c3b73 (
    .a(al_9120ce24),
    .o(al_2ca74a7));
  AL_DFF_1 al_dea139bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2ca74a7),
    .en(1'b1),
    .sr(1'b0),
    .ss(al_b5a5e144),
    .q(al_54b33a69));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    al_8cde73eb (
    .a(al_1e3dbb5f),
    .b(al_bb796872),
    .c(al_5bb559f0),
    .d(al_3f592f2c),
    .o(al_93b093ad[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    al_9af31511 (
    .a(al_b4c6b3bd),
    .b(al_891497d5),
    .c(al_5bb559f0),
    .d(al_3f592f2c),
    .o(al_93b093ad[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    al_3928a88 (
    .a(al_ef78cbcb),
    .b(al_f419b7f2),
    .c(al_5bb559f0),
    .d(al_3f592f2c),
    .o(al_93b093ad[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    al_881cb68b (
    .a(al_d51c2ed1),
    .b(al_f5b9a4c5),
    .c(al_5bb559f0),
    .d(al_3f592f2c),
    .o(al_93b093ad[3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(~D*B)))"),
    .INIT(16'ha028))
    al_36a1a26a (
    .a(al_92b55720[0]),
    .b(al_52b895b5[0]),
    .c(al_52b895b5[1]),
    .d(al_8d73b4c8[0]),
    .o(al_dedaebcb[1]));
  AL_MAP_LUT6 #(
    .EQN("~(E@(~F*D*C*B*A))"),
    .INIT(64'h0000ffff80007fff))
    al_e15a2cdc (
    .a(al_52b895b5[0]),
    .b(al_52b895b5[1]),
    .c(al_52b895b5[2]),
    .d(al_52b895b5[3]),
    .e(al_52b895b5[4]),
    .f(al_8d73b4c8[0]),
    .o(al_fcb84919));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_129acba1 (
    .a(al_fcb84919),
    .b(al_92b55720[0]),
    .o(al_dedaebcb[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_905c81c7 (
    .a(al_fbd177b5),
    .b(al_92b55720[0]),
    .c(al_52b895b5[5]),
    .d(al_52b895b5[6]),
    .e(al_52b895b5[7]),
    .o(al_dedaebcb[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(~D*B)))"),
    .INIT(16'ha028))
    al_88ef2cf (
    .a(al_92b55720[1]),
    .b(al_bd6aead3[0]),
    .c(al_bd6aead3[1]),
    .d(al_8d73b4c8[1]),
    .o(al_6fe26a79[1]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_699017c2 (
    .a(al_47147006),
    .b(al_92b55720[1]),
    .c(al_bd6aead3[2]),
    .d(al_bd6aead3[3]),
    .e(al_bd6aead3[4]),
    .o(al_6fe26a79[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_7013a7f8 (
    .a(al_7b2556ad),
    .b(al_92b55720[1]),
    .c(al_bd6aead3[5]),
    .d(al_bd6aead3[6]),
    .e(al_bd6aead3[7]),
    .o(al_6fe26a79[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(~D*B)))"),
    .INIT(16'ha028))
    al_2f07dfe9 (
    .a(al_92b55720[2]),
    .b(al_febad4d6[0]),
    .c(al_febad4d6[1]),
    .d(al_8d73b4c8[2]),
    .o(al_910cb5e3[1]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_fa119afd (
    .a(al_80311da5),
    .b(al_92b55720[2]),
    .c(al_febad4d6[2]),
    .d(al_febad4d6[3]),
    .e(al_febad4d6[4]),
    .o(al_910cb5e3[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_99b760ed (
    .a(al_c62e8a82),
    .b(al_92b55720[2]),
    .c(al_febad4d6[5]),
    .d(al_febad4d6[6]),
    .e(al_febad4d6[7]),
    .o(al_910cb5e3[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(~D*B)))"),
    .INIT(16'ha028))
    al_4b548c37 (
    .a(al_92b55720[3]),
    .b(al_c57192d3[0]),
    .c(al_c57192d3[1]),
    .d(al_8d73b4c8[3]),
    .o(al_7b9547a0[1]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_8837b636 (
    .a(al_e32a2e7c),
    .b(al_92b55720[3]),
    .c(al_c57192d3[2]),
    .d(al_c57192d3[3]),
    .e(al_c57192d3[4]),
    .o(al_7b9547a0[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_d2bf1d86 (
    .a(al_d31fa142),
    .b(al_92b55720[3]),
    .c(al_c57192d3[5]),
    .d(al_c57192d3[6]),
    .e(al_c57192d3[7]),
    .o(al_7b9547a0[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_4284b0e5 (
    .a(al_92b55720[0]),
    .b(al_52b895b5[0]),
    .c(al_8d73b4c8[0]),
    .o(al_dedaebcb[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_eb9c0f95 (
    .a(al_dedaebcb[5]),
    .b(al_dedaebcb[6]),
    .c(al_dedaebcb[8]),
    .d(al_b6610a70),
    .o(al_e39e8b51[0]));
  AL_MAP_LUT5 #(
    .EQN("(A*(D@(~E*C*B)))"),
    .INIT(32'haa002a80))
    al_a42922df (
    .a(al_92b55720[0]),
    .b(al_52b895b5[0]),
    .c(al_52b895b5[1]),
    .d(al_52b895b5[2]),
    .e(al_8d73b4c8[0]),
    .o(al_dedaebcb[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E@(~F*D*C*B)))"),
    .INIT(64'haaaa00002aaa8000))
    al_c86c3e06 (
    .a(al_92b55720[0]),
    .b(al_52b895b5[0]),
    .c(al_52b895b5[1]),
    .d(al_52b895b5[2]),
    .e(al_52b895b5[3]),
    .f(al_8d73b4c8[0]),
    .o(al_dedaebcb[3]));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*C*B*A)"),
    .INIT(64'h0000000080000000))
    al_cd91ad92 (
    .a(al_52b895b5[0]),
    .b(al_52b895b5[1]),
    .c(al_52b895b5[2]),
    .d(al_52b895b5[3]),
    .e(al_52b895b5[4]),
    .f(al_8d73b4c8[0]),
    .o(al_fbd177b5));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_50a2a911 (
    .a(al_fbd177b5),
    .b(al_92b55720[0]),
    .c(al_52b895b5[5]),
    .o(al_dedaebcb[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_4f42b812 (
    .a(al_fbd177b5),
    .b(al_92b55720[0]),
    .c(al_52b895b5[5]),
    .d(al_52b895b5[6]),
    .o(al_dedaebcb[6]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_d2f6d860 (
    .a(al_fbd177b5),
    .b(al_92b55720[0]),
    .c(al_52b895b5[5]),
    .d(al_52b895b5[6]),
    .e(al_52b895b5[7]),
    .f(al_52b895b5[8]),
    .o(al_dedaebcb[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_cb1888d7 (
    .a(al_dedaebcb[3]),
    .b(al_dedaebcb[2]),
    .c(al_dedaebcb[0]),
    .d(al_52b895b5[1]),
    .e(al_52b895b5[4]),
    .f(al_52b895b5[7]),
    .o(al_b6610a70));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_26918993 (
    .a(al_92b55720[1]),
    .b(al_bd6aead3[0]),
    .c(al_8d73b4c8[1]),
    .o(al_6fe26a79[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_ecb72efc (
    .a(al_1f5470a8),
    .b(al_6fe26a79[5]),
    .c(al_6fe26a79[6]),
    .d(al_6fe26a79[8]),
    .o(al_e39e8b51[1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_f554d808 (
    .a(al_bd6aead3[0]),
    .b(al_bd6aead3[1]),
    .c(al_8d73b4c8[1]),
    .o(al_47147006));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_49ad4efb (
    .a(al_47147006),
    .b(al_92b55720[1]),
    .c(al_bd6aead3[2]),
    .o(al_6fe26a79[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_28c75f11 (
    .a(al_47147006),
    .b(al_92b55720[1]),
    .c(al_bd6aead3[2]),
    .d(al_bd6aead3[3]),
    .o(al_6fe26a79[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_cb179044 (
    .a(al_47147006),
    .b(al_bd6aead3[2]),
    .c(al_bd6aead3[3]),
    .d(al_bd6aead3[4]),
    .o(al_7b2556ad));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_bf13f61 (
    .a(al_7b2556ad),
    .b(al_92b55720[1]),
    .c(al_bd6aead3[5]),
    .o(al_6fe26a79[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_59365ca6 (
    .a(al_7b2556ad),
    .b(al_92b55720[1]),
    .c(al_bd6aead3[5]),
    .d(al_bd6aead3[6]),
    .o(al_6fe26a79[6]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_53f2411d (
    .a(al_7b2556ad),
    .b(al_92b55720[1]),
    .c(al_bd6aead3[5]),
    .d(al_bd6aead3[6]),
    .e(al_bd6aead3[7]),
    .f(al_bd6aead3[8]),
    .o(al_6fe26a79[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_83f43007 (
    .a(al_6fe26a79[2]),
    .b(al_6fe26a79[3]),
    .c(al_6fe26a79[0]),
    .d(al_bd6aead3[1]),
    .e(al_bd6aead3[4]),
    .f(al_bd6aead3[7]),
    .o(al_1f5470a8));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_bdd6be1c (
    .a(al_92b55720[2]),
    .b(al_febad4d6[0]),
    .c(al_8d73b4c8[2]),
    .o(al_910cb5e3[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_ee20a233 (
    .a(al_f100fb27),
    .b(al_910cb5e3[5]),
    .c(al_910cb5e3[6]),
    .d(al_910cb5e3[8]),
    .o(al_e39e8b51[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_90957ef9 (
    .a(al_febad4d6[0]),
    .b(al_febad4d6[1]),
    .c(al_8d73b4c8[2]),
    .o(al_80311da5));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_8a31c4a2 (
    .a(al_80311da5),
    .b(al_92b55720[2]),
    .c(al_febad4d6[2]),
    .o(al_910cb5e3[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_c6620303 (
    .a(al_80311da5),
    .b(al_92b55720[2]),
    .c(al_febad4d6[2]),
    .d(al_febad4d6[3]),
    .o(al_910cb5e3[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_81f20fed (
    .a(al_80311da5),
    .b(al_febad4d6[2]),
    .c(al_febad4d6[3]),
    .d(al_febad4d6[4]),
    .o(al_c62e8a82));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_5fa98ab2 (
    .a(al_c62e8a82),
    .b(al_92b55720[2]),
    .c(al_febad4d6[5]),
    .o(al_910cb5e3[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_69a660e5 (
    .a(al_c62e8a82),
    .b(al_92b55720[2]),
    .c(al_febad4d6[5]),
    .d(al_febad4d6[6]),
    .o(al_910cb5e3[6]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_42be2206 (
    .a(al_c62e8a82),
    .b(al_92b55720[2]),
    .c(al_febad4d6[5]),
    .d(al_febad4d6[6]),
    .e(al_febad4d6[7]),
    .f(al_febad4d6[8]),
    .o(al_910cb5e3[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_59d23c63 (
    .a(al_910cb5e3[2]),
    .b(al_910cb5e3[3]),
    .c(al_910cb5e3[0]),
    .d(al_febad4d6[1]),
    .e(al_febad4d6[4]),
    .f(al_febad4d6[7]),
    .o(al_f100fb27));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_9b634b3a (
    .a(al_92b55720[3]),
    .b(al_c57192d3[0]),
    .c(al_8d73b4c8[3]),
    .o(al_7b9547a0[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_deb3e38c (
    .a(al_ac3a915e),
    .b(al_7b9547a0[5]),
    .c(al_7b9547a0[6]),
    .d(al_7b9547a0[8]),
    .o(al_e39e8b51[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_caf2bcba (
    .a(al_c57192d3[0]),
    .b(al_c57192d3[1]),
    .c(al_8d73b4c8[3]),
    .o(al_e32a2e7c));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_7d7afa1 (
    .a(al_e32a2e7c),
    .b(al_92b55720[3]),
    .c(al_c57192d3[2]),
    .o(al_7b9547a0[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_c612fe1f (
    .a(al_e32a2e7c),
    .b(al_92b55720[3]),
    .c(al_c57192d3[2]),
    .d(al_c57192d3[3]),
    .o(al_7b9547a0[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_3a9ca0af (
    .a(al_e32a2e7c),
    .b(al_c57192d3[2]),
    .c(al_c57192d3[3]),
    .d(al_c57192d3[4]),
    .o(al_d31fa142));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_5286705 (
    .a(al_d31fa142),
    .b(al_92b55720[3]),
    .c(al_c57192d3[5]),
    .o(al_7b9547a0[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_14fab9a8 (
    .a(al_d31fa142),
    .b(al_92b55720[3]),
    .c(al_c57192d3[5]),
    .d(al_c57192d3[6]),
    .o(al_7b9547a0[6]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_ee84ed0c (
    .a(al_d31fa142),
    .b(al_92b55720[3]),
    .c(al_c57192d3[5]),
    .d(al_c57192d3[6]),
    .e(al_c57192d3[7]),
    .f(al_c57192d3[8]),
    .o(al_7b9547a0[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_d9fb74ce (
    .a(al_7b9547a0[2]),
    .b(al_7b9547a0[3]),
    .c(al_7b9547a0[0]),
    .d(al_c57192d3[1]),
    .e(al_c57192d3[4]),
    .f(al_c57192d3[7]),
    .o(al_ac3a915e));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_6d04d850 (
    .a(al_b5a5e144),
    .b(al_ef9accde),
    .c(al_6ad27cba[0]),
    .d(al_6ad27cba[1]),
    .o(al_6a03de0));
  AL_DFF_0 al_ea983e44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6a03de0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6ad27cba[0]));
  AL_DFF_0 al_345ec426 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_efc928b8[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_6ad27cba[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_33fe61f6 (
    .a(al_ef9accde),
    .b(al_6ad27cba[1]),
    .o(al_99917cb7));
  AL_DFF_1 al_717b9ebc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_99917cb7),
    .en(1'b1),
    .sr(1'b0),
    .ss(al_b5a5e144),
    .q(al_c9d121b2));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    al_a72ca3ff (
    .a(al_ef9accde),
    .b(al_6ad27cba[0]),
    .c(al_6ad27cba[1]),
    .o(al_efc928b8[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_a43dcbe (
    .a(al_90b7699),
    .b(al_c58e2364[0]),
    .o(al_97b2c696[0]));
  AL_MAP_LUT5 #(
    .EQN("~(~D*C*A*~(~E*B))"),
    .INIT(32'hff5fffdf))
    al_b208e581 (
    .a(al_9941dfb9[0]),
    .b(al_9941dfb9[1]),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .e(al_c5fa5405),
    .o(al_c18a6fab));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A*~(D@C)))"),
    .INIT(16'hb33b))
    al_1bd2c570 (
    .a(al_8e57b8ea),
    .b(al_c18a6fab),
    .c(al_c58e2364[0]),
    .d(al_c58e2364[1]),
    .o(al_97b2c696[1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(~C*~B)))"),
    .INIT(16'ha802))
    al_51df63b3 (
    .a(al_90b7699),
    .b(al_c58e2364[0]),
    .c(al_c58e2364[1]),
    .d(al_c58e2364[2]),
    .o(al_97b2c696[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_34bc9d47 (
    .a(al_bc505469[0]),
    .b(al_bc505469[1]),
    .c(al_bc505469[2]),
    .d(al_bc505469[3]),
    .o(al_cb6618b2));
  AL_MAP_LUT5 #(
    .EQN("(~A*(~(B)*~(C)*~(D)*~(E)+B*~(C)*~(D)*~(E)+~(B)*C*~(D)*~(E)+~(B)*C*D*~(E)+B*C*D*~(E)+B*~(C)*~(D)*E+~(B)*C*~(D)*E+~(B)*~(C)*D*E+B*~(C)*D*E+~(B)*C*D*E+B*C*D*E))"),
    .INIT(32'h55145015))
    al_e9440f9 (
    .a(al_eb540174),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .o(al_8e57b8ea));
  AL_MAP_LUT6 #(
    .EQN("(~E*D*B*(~A*~(F)*~(C)+~A*F*~(C)+~(~A)*F*C+~A*F*C))"),
    .INIT(64'h0000c40000000400))
    al_76955a88 (
    .a(al_cb6618b2),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_c5fa5405),
    .o(al_3225efe4));
  AL_MAP_LUT6 #(
    .EQN("~(~B*~(A*(F@(~E*~D*~C))))"),
    .INIT(64'heeeeeeecccccccce))
    al_f9e7f9fa (
    .a(al_8e57b8ea),
    .b(al_3225efe4),
    .c(al_c58e2364[0]),
    .d(al_c58e2364[1]),
    .e(al_c58e2364[2]),
    .f(al_c58e2364[3]),
    .o(al_97b2c696[3]));
  AL_MAP_LUT6 #(
    .EQN("(~A*(F@(~E*~D*~C*~B)))"),
    .INIT(64'h5555555400000001))
    al_e35ce9be (
    .a(al_eb540174),
    .b(al_c58e2364[0]),
    .c(al_c58e2364[1]),
    .d(al_c58e2364[2]),
    .e(al_c58e2364[3]),
    .f(al_c58e2364[4]),
    .o(al_18ebfba6));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haaeb2c2aaaebac2a))
    al_b006c13a (
    .a(al_18ebfba6),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_c5fa5405),
    .o(al_97b2c696[4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_64002775 (
    .a(al_2d8af247),
    .b(al_c58e2364[5]),
    .c(al_c58e2364[6]),
    .d(al_c58e2364[7]),
    .o(al_eb540174));
  AL_MAP_LUT6 #(
    .EQN("(~A*(~(B)*~(C)*~(D)*~(E)*~(F)+B*~(C)*~(D)*~(E)*~(F)+~(B)*C*~(D)*~(E)*~(F)+~(B)*C*D*~(E)*~(F)+B*C*D*~(E)*~(F)+B*~(C)*~(D)*E*~(F)+~(B)*C*~(D)*E*~(F)+~(B)*~(C)*D*E*~(F)+B*~(C)*D*E*~(F)+~(B)*C*D*E*~(F)+B*C*D*E*~(F)+~(B)*~(C)*~(D)*~(E)*F+B*~(C)*~(D)*~(E)*F+~(B)*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*~(C)*~(D)*E*F+~(B)*C*~(D)*E*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'h5514101555145015))
    al_f2f4d481 (
    .a(al_eb540174),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_c5fa5405),
    .o(al_90b7699));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    al_c633b5e7 (
    .a(al_90b7699),
    .b(al_2d8af247),
    .c(al_c58e2364[5]),
    .o(al_97b2c696[5]));
  AL_MAP_LUT4 #(
    .EQN("(~((~B*A))*~(C)*~(D)+(~B*A)*~(C)*~(D)+(~B*A)*C*~(D)+~((~B*A))*~(C)*D+(~B*A)*C*D)"),
    .INIT(16'h2d2f))
    al_7c68c855 (
    .a(al_2d8af247),
    .b(al_c58e2364[5]),
    .c(al_c58e2364[6]),
    .d(al_c58e2364[7]),
    .o(al_e3c7998c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h55d4101555d45015))
    al_b41f22ee (
    .a(al_e3c7998c),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_c5fa5405),
    .o(al_97b2c696[6]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_f2d64b9 (
    .a(al_c58e2364[0]),
    .b(al_c58e2364[1]),
    .c(al_c58e2364[2]),
    .d(al_c58e2364[3]),
    .e(al_c58e2364[4]),
    .o(al_2d8af247));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    al_81d634d2 (
    .a(al_2d8af247),
    .b(al_c58e2364[5]),
    .c(al_c58e2364[6]),
    .d(al_c58e2364[7]),
    .o(al_c7a09c4f));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haae8202aaae8a02a))
    al_5b6e93c4 (
    .a(al_c7a09c4f),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_c5fa5405),
    .o(al_97b2c696[7]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*D*C*B))"),
    .INIT(32'h2aaaaaaa))
    al_810a9b08 (
    .a(al_3bfb3478),
    .b(al_2f365000[0]),
    .c(al_2f365000[1]),
    .d(al_2f365000[2]),
    .e(al_2f365000[3]),
    .o(al_72e5ab2f));
  AL_DFF_0 al_35052a43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_72e5ab2f),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_d9786abc));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*~B*~A)"),
    .INIT(32'h00000100))
    al_35f1ddac (
    .a(al_b5a5e144),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .o(al_8514591d));
  AL_DFF_0 al_1c1e825c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8514591d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f7a36e8));
  AL_DFF_0 al_f408ed80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9821c430),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c5705f8a));
  AL_MAP_LUT6 #(
    .EQN("(~B*~A*~(~F*~E*~D*~C))"),
    .INIT(64'h1111111111111110))
    al_341bf8fe (
    .a(al_cf11b78b[2]),
    .b(al_a082bc48),
    .c(al_2f365000[0]),
    .d(al_2f365000[1]),
    .e(al_2f365000[2]),
    .f(al_2f365000[3]),
    .o(al_62d3bb1d));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_de7d4da0 (
    .a(al_62d3bb1d),
    .b(al_cf11b78b[0]),
    .c(al_cf11b78b[1]),
    .d(al_cf11b78b[3]),
    .o(al_21374d40));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hcccc0cccc0cccecc))
    al_9d21685 (
    .a(al_21374d40),
    .b(al_898823b1),
    .c(al_9941dfb9[0]),
    .d(al_9941dfb9[1]),
    .e(al_9941dfb9[2]),
    .f(al_9941dfb9[3]),
    .o(al_731b9711));
  AL_DFF_0 al_e3ec0aee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_731b9711),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_898823b1));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~((F*~E))+A*B*~(C)*~(D)*~((F*~E))+~(A)*B*C*~(D)*~((F*~E))+A*B*C*~(D)*~((F*~E))+~(A)*B*~(C)*D*~((F*~E))+A*B*~(C)*D*~((F*~E))+~(A)*B*C*D*~((F*~E))+A*B*C*D*~((F*~E))+~(A)*B*~(C)*~(D)*(F*~E)+A*B*~(C)*~(D)*(F*~E)+~(A)*~(B)*C*~(D)*(F*~E)+A*~(B)*C*~(D)*(F*~E)+~(A)*B*C*~(D)*(F*~E)+A*B*C*~(D)*(F*~E)+A*B*~(C)*D*(F*~E))"),
    .INIT(64'hcccc08fccccccccc))
    al_ca8e5a6a (
    .a(init_calib_complete),
    .b(al_79090ab6),
    .c(al_9941dfb9[0]),
    .d(al_9941dfb9[1]),
    .e(al_9941dfb9[2]),
    .f(al_9941dfb9[3]),
    .o(al_1cd23aa7));
  AL_DFF_0 al_36c245e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1cd23aa7),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_79090ab6));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*~A)"),
    .INIT(32'h00400000))
    al_e51f96d2 (
    .a(al_b5a5e144),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .o(al_c1a95cc7));
  AL_DFF_0 al_67b4f0d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c1a95cc7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41c9267e));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    al_1e6340cc (
    .a(al_b5a5e144),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .o(al_4566fdd3));
  AL_DFF_0 al_dad92f10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4566fdd3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11b28491));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*C*~D+A*B*~C*D)"),
    .INIT(16'b0000100000100000))
    al_a6616b1b (
    .a(al_9941dfb9[0]),
    .b(al_9941dfb9[1]),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .o(al_9821c430));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_69e2df84 (
    .a(al_aca36a53),
    .b(al_b5a5e144),
    .o(al_49733697));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E@(~(B)*C*~(D)+B*~(C)*D)))"),
    .INIT(32'hfbefaeba))
    al_df39b7ed (
    .a(al_4bd4fa38),
    .b(al_d9786abc),
    .c(al_4f7a36e8),
    .d(al_2f365000[0]),
    .e(al_2f365000[1]),
    .o(al_c9543684[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(C)*~(D)*~((~E*B))+A*~(C)*~(D)*~((~E*B))+~(A)*~(C)*D*~((~E*B))+~(A)*~(C)*~(D)*(~E*B)+A*~(C)*~(D)*(~E*B)+~(A)*C*~(D)*(~E*B)+A*C*~(D)*(~E*B)+~(A)*~(C)*D*(~E*B))"),
    .INIT(32'h050f05cf))
    al_1d7e3771 (
    .a(al_21374d40),
    .b(al_eb540174),
    .c(al_9941dfb9[0]),
    .d(al_9941dfb9[1]),
    .e(al_a769a364[0]),
    .o(al_ac57883f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffc3cf55ffc30f55))
    al_9447e723 (
    .a(al_ac57883f),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_c5fa5405),
    .o(al_b4db00cd[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_e5f4e457 (
    .a(al_cf11b78b[0]),
    .b(al_cf11b78b[1]),
    .c(al_cf11b78b[2]),
    .d(al_cf11b78b[3]),
    .o(al_28570942));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*C*~(D)*~(E)*~((F*A))+B*C*~(D)*~(E)*~((F*A))+~(B)*~(C)*~(D)*E*~((F*A))+B*~(C)*~(D)*E*~((F*A))+~(B)*C*~(D)*E*~((F*A))+B*C*~(D)*E*~((F*A))+~(B)*~(C)*D*E*~((F*A))+~(B)*C*D*E*~((F*A))+~(B)*C*~(D)*~(E)*(F*A)+B*C*~(D)*~(E)*(F*A)+~(B)*~(C)*D*~(E)*(F*A)+B*~(C)*D*~(E)*(F*A)+~(B)*C*D*~(E)*(F*A)+B*C*D*~(E)*(F*A)+~(B)*~(C)*~(D)*E*(F*A)+B*~(C)*~(D)*E*(F*A)+~(B)*C*~(D)*E*(F*A)+B*C*~(D)*E*(F*A)+~(B)*~(C)*D*E*(F*A)+~(B)*C*D*E*(F*A))"),
    .INIT(64'h33ffaaf033ff00f0))
    al_c334fe5a (
    .a(al_eb540174),
    .b(al_28570942),
    .c(init_calib_complete),
    .d(al_9941dfb9[0]),
    .e(al_9941dfb9[1]),
    .f(al_a769a364[1]),
    .o(al_cc80b352));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00d3cfff00d30fff))
    al_313f35a1 (
    .a(init_calib_complete),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_c5fa5405),
    .o(al_4e9593a4));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(~D*~C*A))"),
    .INIT(16'h333b))
    al_d10457d9 (
    .a(al_cc80b352),
    .b(al_4e9593a4),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .o(al_b4db00cd[1]));
  AL_MAP_LUT6 #(
    .EQN("~(B*(C*D*~((E*A))*~(F)+~(C)*~(D)*(E*A)*~(F)+C*D*(E*A)*~(F)+~(C)*~(D)*(E*A)*F))"),
    .INIT(64'hfff7ffff3ff73fff))
    al_ec057a7e (
    .a(al_eb540174),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_a769a364[2]),
    .f(al_c5fa5405),
    .o(al_7941134));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_4beb6f37 (
    .a(al_7941134),
    .b(al_9941dfb9[2]),
    .c(al_9941dfb9[3]),
    .o(al_b4db00cd[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_d8677c9d (
    .a(al_eb540174),
    .b(al_9941dfb9[2]),
    .c(al_9941dfb9[3]),
    .d(al_a769a364[3]),
    .o(al_a6b572a3));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffff0cf000a000a0))
    al_2181ade4 (
    .a(al_a6b572a3),
    .b(init_calib_complete),
    .c(al_9941dfb9[0]),
    .d(al_9941dfb9[1]),
    .e(al_9941dfb9[2]),
    .f(al_9941dfb9[3]),
    .o(al_b4db00cd[3]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C@B))"),
    .INIT(8'hbe))
    al_fb7da254 (
    .a(al_3bfb3478),
    .b(init_calib_complete),
    .c(al_48a3872d[0]),
    .o(al_55d92da7[0]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D@(~C*B)))"),
    .INIT(16'hfbae))
    al_1f10f3c6 (
    .a(al_3bfb3478),
    .b(init_calib_complete),
    .c(al_48a3872d[0]),
    .d(al_48a3872d[1]),
    .o(al_55d92da7[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(E@(~D*~C*B)))"),
    .INIT(32'h55510004))
    al_82077ad5 (
    .a(al_3bfb3478),
    .b(init_calib_complete),
    .c(al_48a3872d[0]),
    .d(al_48a3872d[1]),
    .e(al_48a3872d[2]),
    .o(al_55d92da7[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffdf0830))
    al_3ea1850b (
    .a(al_9941dfb9[0]),
    .b(al_9941dfb9[1]),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .e(al_bc505469[0]),
    .o(al_df310708[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf7eff7cf00000020))
    al_968cc5b0 (
    .a(al_9941dfb9[0]),
    .b(al_9941dfb9[1]),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .e(al_bc505469[0]),
    .f(al_bc505469[1]),
    .o(al_df310708[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3ff4ff00000800))
    al_550c6117 (
    .a(al_3e848d66),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_bc505469[2]),
    .o(al_df310708[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_fcf19fc3 (
    .a(al_bc505469[0]),
    .b(al_bc505469[1]),
    .o(al_3e848d66));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_834b025f (
    .a(al_3e848d66),
    .b(al_bc505469[2]),
    .o(al_42f2763a));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3ff4ff00000800))
    al_1846e8d3 (
    .a(al_42f2763a),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_bc505469[3]),
    .o(al_df310708[3]));
  AL_DFF_1 al_bd4164b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[0]));
  AL_DFF_1 al_f295f5f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[1]));
  AL_DFF_1 al_3aced2fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[2]));
  AL_DFF_1 al_a25f1b8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[3]));
  AL_DFF_1 al_ff09ce21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[4]));
  AL_DFF_1 al_74bbfb93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[5]));
  AL_DFF_1 al_3457d0c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[6]));
  AL_DFF_1 al_a108f1f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[7]));
  AL_DFF_1 al_e3401ea9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[8]));
  AL_DFF_1 al_6a7ccd00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[9]));
  AL_DFF_1 al_4b964d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[10]));
  AL_DFF_1 al_b05850e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[11]));
  AL_DFF_1 al_37ae219 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[12]));
  AL_DFF_1 al_20b77a84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[13]));
  AL_DFF_1 al_b4132867 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[14]));
  AL_DFF_1 al_b636370c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a27c86[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(~al_49733697),
    .q(al_e827ceba[15]));
  AL_DFF_0 al_4b9fa95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97b2c696[0]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58e2364[0]));
  AL_DFF_0 al_d9c8c824 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97b2c696[1]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58e2364[1]));
  AL_DFF_0 al_593340 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97b2c696[2]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58e2364[2]));
  AL_DFF_0 al_44d4cebe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97b2c696[3]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58e2364[3]));
  AL_DFF_0 al_99369454 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97b2c696[4]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58e2364[4]));
  AL_DFF_0 al_2de7826b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97b2c696[5]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58e2364[5]));
  AL_DFF_0 al_ed67a6c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97b2c696[6]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58e2364[6]));
  AL_DFF_0 al_a0bcfa97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_97b2c696[7]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c58e2364[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_af168aa2 (
    .a(al_d9786abc),
    .b(al_2f365000[0]),
    .c(al_2f365000[1]),
    .o(al_d0f70b25[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*(~(A)*~(C)*~(D)+A*C*D))"),
    .INIT(16'h8004))
    al_dd4a323d (
    .a(al_d9786abc),
    .b(al_4f7a36e8),
    .c(al_2f365000[0]),
    .d(al_2f365000[1]),
    .o(al_ad018368));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*(B@A))"),
    .INIT(16'h0600))
    al_f32b96a6 (
    .a(al_9941dfb9[0]),
    .b(al_9941dfb9[1]),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .o(al_4bd4fa38));
  AL_MAP_LUT5 #(
    .EQN("(~B*~A*(E@D@C))"),
    .INIT(32'h10010110))
    al_6bd0fc95 (
    .a(al_4bd4fa38),
    .b(al_b5a5e144),
    .c(al_d9786abc),
    .d(al_4f7a36e8),
    .e(al_2f365000[0]),
    .o(al_2957c84b));
  AL_MAP_LUT5 #(
    .EQN("(~D*~B*(E@C@A))"),
    .INIT(32'h00210012))
    al_91c2b295 (
    .a(al_ad018368),
    .b(al_4bd4fa38),
    .c(al_d0f70b25[1]),
    .d(al_b5a5e144),
    .e(al_2f365000[2]),
    .o(al_c79b855c));
  AL_MAP_LUT6 #(
    .EQN("(~D*~B*(F@(A*~(C)*~(E)+~(A)*C*E)))"),
    .INIT(64'h0023003100100002))
    al_c6080bc2 (
    .a(al_ad018368),
    .b(al_4bd4fa38),
    .c(al_d0f70b25[1]),
    .d(al_b5a5e144),
    .e(al_2f365000[2]),
    .f(al_2f365000[3]),
    .o(al_3ac9505a));
  AL_DFF_0 al_9ac8b07a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2957c84b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f365000[0]));
  AL_DFF_0 al_89233af5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c9543684[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_2f365000[1]));
  AL_DFF_0 al_55d6c675 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c79b855c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f365000[2]));
  AL_DFF_0 al_db0c06ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3ac9505a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f365000[3]));
  AL_DFF_0 al_a3650c2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4db00cd[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_9941dfb9[0]));
  AL_DFF_0 al_4b451c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4db00cd[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_9941dfb9[1]));
  AL_DFF_0 al_4afbc6a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4db00cd[2]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_9941dfb9[2]));
  AL_DFF_0 al_415b03ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4db00cd[3]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_9941dfb9[3]));
  AL_DFF_0 al_847d8ba6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55d92da7[0]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_48a3872d[0]));
  AL_DFF_0 al_e396f7da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55d92da7[1]),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_48a3872d[1]));
  AL_DFF_0 al_8e5aa8d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_434e6eb1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48a3872d[4]));
  AL_DFF_0 al_7030ad25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_365f3d23),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48a3872d[5]));
  AL_DFF_0 al_2a317c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0784ca8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48a3872d[6]));
  AL_DFF_0 al_578c71de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_badd7923),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48a3872d[7]));
  AL_DFF_1 al_6aaedb00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55d92da7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(al_b5a5e144),
    .q(al_48a3872d[2]));
  AL_DFF_1 al_92b28b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_79c695eb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48a3872d[3]));
  AL_DFF_1 al_a0293694 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3a7e0263),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48a3872d[8]));
  AL_DFF_1 al_b43d83dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9a44af5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48a3872d[9]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_7da198e3 (
    .a(al_48a3872d[0]),
    .b(al_48a3872d[1]),
    .c(al_48a3872d[4]),
    .d(al_48a3872d[5]),
    .e(al_48a3872d[6]),
    .f(al_48a3872d[7]),
    .o(al_4ae2fdc2));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_78405df4 (
    .a(al_4ae2fdc2),
    .b(al_48a3872d[2]),
    .c(al_48a3872d[3]),
    .d(al_48a3872d[8]),
    .e(al_48a3872d[9]),
    .o(al_3bfb3478));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_d52a0313 (
    .a(init_calib_complete),
    .b(al_48a3872d[0]),
    .c(al_48a3872d[1]),
    .d(al_48a3872d[4]),
    .e(al_48a3872d[2]),
    .f(al_48a3872d[3]),
    .o(al_9b29508b));
  AL_MAP_LUT6 #(
    .EQN("~(D@(~F*~E*~C*~B*A))"),
    .INIT(64'h00ff00ff00ff02fd))
    al_538c0009 (
    .a(init_calib_complete),
    .b(al_48a3872d[0]),
    .c(al_48a3872d[1]),
    .d(al_48a3872d[4]),
    .e(al_48a3872d[2]),
    .f(al_48a3872d[3]),
    .o(al_db03633e));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_4546c08c (
    .a(al_3bfb3478),
    .b(al_b5a5e144),
    .o(al_fe37e390));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_72ea90a7 (
    .a(al_fe37e390),
    .b(al_db03633e),
    .o(al_434e6eb1));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    al_c77d0df1 (
    .a(al_fe37e390),
    .b(al_9b29508b),
    .c(al_48a3872d[5]),
    .o(al_365f3d23));
  AL_MAP_LUT6 #(
    .EQN("~(A*~(F@(~E*~D*~C*B)))"),
    .INIT(64'hfffffff75555555d))
    al_f215be7b (
    .a(al_fe37e390),
    .b(init_calib_complete),
    .c(al_48a3872d[0]),
    .d(al_48a3872d[1]),
    .e(al_48a3872d[2]),
    .f(al_48a3872d[3]),
    .o(al_79c695eb));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(~C*B)))"),
    .INIT(16'ha208))
    al_fc5b2c2d (
    .a(al_fe37e390),
    .b(al_9b29508b),
    .c(al_48a3872d[5]),
    .d(al_48a3872d[6]),
    .o(al_b0784ca8));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@(~D*~C*B)))"),
    .INIT(32'haaa20008))
    al_f9ef9fa4 (
    .a(al_fe37e390),
    .b(al_9b29508b),
    .c(al_48a3872d[5]),
    .d(al_48a3872d[6]),
    .e(al_48a3872d[7]),
    .o(al_badd7923));
  AL_MAP_LUT6 #(
    .EQN("~(A*~(F@(~E*~D*~C*B)))"),
    .INIT(64'hfffffff75555555d))
    al_c0654183 (
    .a(al_fe37e390),
    .b(al_9b29508b),
    .c(al_48a3872d[5]),
    .d(al_48a3872d[6]),
    .e(al_48a3872d[7]),
    .f(al_48a3872d[8]),
    .o(al_3a7e0263));
  AL_MAP_LUT6 #(
    .EQN("(F@(~E*~D*~C*~B*A))"),
    .INIT(64'hfffffffd00000002))
    al_37dd8c3 (
    .a(al_9b29508b),
    .b(al_48a3872d[5]),
    .c(al_48a3872d[6]),
    .d(al_48a3872d[7]),
    .e(al_48a3872d[8]),
    .f(al_48a3872d[9]),
    .o(al_a923bd8[9]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    al_6f4a4707 (
    .a(al_fe37e390),
    .b(al_a923bd8[9]),
    .o(al_9a44af5));
  AL_DFF_0 al_3063117c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_df310708[0]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bc505469[0]));
  AL_DFF_0 al_4768a0e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_df310708[1]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bc505469[1]));
  AL_DFF_0 al_e1d852f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_df310708[2]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bc505469[2]));
  AL_DFF_0 al_6bbe54ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_df310708[3]),
    .en(al_9388375e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bc505469[3]));
  AL_DFF_0 al_8e7a22d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b4486c6[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a769a364[0]));
  AL_DFF_0 al_4ac40b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b4486c6[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a769a364[1]));
  AL_DFF_0 al_a79fe38a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b4486c6[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a769a364[2]));
  AL_DFF_0 al_d08623f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b4486c6[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a769a364[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfe770830fef70830))
    al_6b251325 (
    .a(al_9941dfb9[0]),
    .b(al_9941dfb9[1]),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .e(al_a769a364[0]),
    .f(al_c5fa5405),
    .o(al_8b4486c6[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc7f707f7))
    al_7db29dc5 (
    .a(al_cb6618b2),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_a769a364[1]),
    .e(al_c5fa5405),
    .o(al_fff872b2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3f553f00035500))
    al_f5a5e11d (
    .a(al_fff872b2),
    .b(al_9941dfb9[0]),
    .c(al_9941dfb9[1]),
    .d(al_9941dfb9[2]),
    .e(al_9941dfb9[3]),
    .f(al_a769a364[1]),
    .o(al_8b4486c6[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff7f0938ffff0938))
    al_518ca330 (
    .a(al_9941dfb9[0]),
    .b(al_9941dfb9[1]),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .e(al_a769a364[2]),
    .f(al_c5fa5405),
    .o(al_8b4486c6[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf6c70080f6c70000))
    al_a220126 (
    .a(al_9941dfb9[0]),
    .b(al_9941dfb9[1]),
    .c(al_9941dfb9[2]),
    .d(al_9941dfb9[3]),
    .e(al_a769a364[3]),
    .f(al_c5fa5405),
    .o(al_8b4486c6[3]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_4f65094c (
    .a(1'b0),
    .o({al_743fb5ed,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cf0f6b01 (
    .a(al_e827ceba[0]),
    .b(al_c5705f8a),
    .c(al_743fb5ed),
    .o({al_c8295b95,al_4a27c86[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_88b52457 (
    .a(al_e827ceba[1]),
    .b(1'b0),
    .c(al_c8295b95),
    .o({al_ec4a81f,al_4a27c86[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c8efedb1 (
    .a(al_e827ceba[2]),
    .b(1'b0),
    .c(al_ec4a81f),
    .o({al_40d806bd,al_4a27c86[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbfab65f (
    .a(al_e827ceba[3]),
    .b(1'b0),
    .c(al_40d806bd),
    .o({al_45a34621,al_4a27c86[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a8cbcb0a (
    .a(al_e827ceba[4]),
    .b(1'b0),
    .c(al_45a34621),
    .o({al_cb5fd325,al_4a27c86[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_365e2688 (
    .a(al_e827ceba[5]),
    .b(1'b0),
    .c(al_cb5fd325),
    .o({al_9680139f,al_4a27c86[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_344fbd88 (
    .a(al_e827ceba[6]),
    .b(1'b0),
    .c(al_9680139f),
    .o({al_7d50905e,al_4a27c86[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a7f2a3 (
    .a(al_e827ceba[7]),
    .b(1'b0),
    .c(al_7d50905e),
    .o({al_92e38148,al_4a27c86[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b3e5c805 (
    .a(al_e827ceba[8]),
    .b(1'b0),
    .c(al_92e38148),
    .o({al_eb5035c8,al_4a27c86[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6f6222ca (
    .a(al_e827ceba[9]),
    .b(1'b0),
    .c(al_eb5035c8),
    .o({al_6cc9e68d,al_4a27c86[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_80bf313 (
    .a(al_e827ceba[10]),
    .b(1'b0),
    .c(al_6cc9e68d),
    .o({al_ca0e45f8,al_4a27c86[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d02d1a27 (
    .a(al_e827ceba[11]),
    .b(1'b0),
    .c(al_ca0e45f8),
    .o({al_f44df3e,al_4a27c86[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a336cb1a (
    .a(al_e827ceba[12]),
    .b(1'b0),
    .c(al_f44df3e),
    .o({al_d7181d37,al_4a27c86[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_805c81b (
    .a(al_e827ceba[13]),
    .b(1'b0),
    .c(al_d7181d37),
    .o({al_c3029dcc,al_4a27c86[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_82ea7554 (
    .a(al_e827ceba[14]),
    .b(1'b0),
    .c(al_c3029dcc),
    .o({al_3ba0cc79,al_4a27c86[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_21798b66 (
    .a(al_e827ceba[15]),
    .b(1'b0),
    .c(al_3ba0cc79),
    .o({open_n11,al_4a27c86[15]}));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_3e9bd74e (
    .a(al_e827ceba[0]),
    .b(al_e827ceba[1]),
    .c(al_e827ceba[2]),
    .d(al_e827ceba[3]),
    .o(al_acfaa45c));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_bb27fe24 (
    .a(al_e827ceba[8]),
    .b(al_e827ceba[9]),
    .c(al_e827ceba[10]),
    .d(al_e827ceba[11]),
    .o(al_a83cb045));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_af792581 (
    .a(al_a83cb045),
    .b(al_e827ceba[12]),
    .c(al_e827ceba[13]),
    .d(al_e827ceba[14]),
    .e(al_e827ceba[15]),
    .o(al_c1f0ed98));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_30201442 (
    .a(al_c1f0ed98),
    .b(al_acfaa45c),
    .c(al_e827ceba[4]),
    .d(al_e827ceba[5]),
    .e(al_e827ceba[6]),
    .f(al_e827ceba[7]),
    .o(al_aca36a53));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    al_9c3dcf78 (
    .a(al_aca36a53),
    .b(al_11b28491),
    .c(al_c5fa5405),
    .o(al_dcd8888a));
  AL_DFF_0 al_f7c646d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dcd8888a),
    .en(1'b1),
    .sr(al_b5a5e144),
    .ss(1'b0),
    .q(al_c5fa5405));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a36b55ba (
    .i(al_a3c26eaf),
    .o(al_813c693b));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_8df72a60 (
    .i(al_813c693b),
    .o(al_6db5b9d2));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_b07d861a (
    .a(ddr_app_en),
    .b(ddr_app_rdy),
    .o(al_e58efc01));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT(16'h2230))
    al_9115b5a8 (
    .a(ddr_app_en),
    .b(al_6db5b9d2),
    .c(al_489041e9),
    .d(ddr_app_rdy),
    .o(al_bf594241));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h4450))
    al_84a5b9ac (
    .a(al_6db5b9d2),
    .b(al_489041e9),
    .c(al_61f44420),
    .d(ddr_app_rdy),
    .o(al_10f4d190));
  AL_DFF_0 al_2161dfd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bf594241),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_489041e9));
  AL_DFF_0 al_97e177f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_10f4d190),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_61f44420));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_17de0460 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[3]),
    .c(al_5d3f410a[3]),
    .o(al_58fb4752[3]));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(~C*A))"),
    .INIT(16'h39c6))
    al_14ee6c19 (
    .a(al_864a13d9[0]),
    .b(al_864a13d9[1]),
    .c(al_f2dedfad[0]),
    .d(al_f2dedfad[1]),
    .o(al_54004a97));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*~B*~A)"),
    .INIT(32'h00001000))
    al_6a0f1485 (
    .a(al_54004a97),
    .b(al_58fb4752[3]),
    .c(al_58fb4752[4]),
    .d(init_calib_complete),
    .e(al_7c9229ee),
    .o(al_40276cd4));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(~C*A))"),
    .INIT(16'h39c6))
    al_acf1fa2b (
    .a(al_b1a73cf[0]),
    .b(al_b1a73cf[1]),
    .c(al_1124d2df[0]),
    .d(al_1124d2df[1]),
    .o(al_5a6db454));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*~A)"),
    .INIT(32'h00004000))
    al_a0e6c5a5 (
    .a(al_5a6db454),
    .b(al_58fb4752[3]),
    .c(al_58fb4752[4]),
    .d(init_calib_complete),
    .e(al_7c9229ee),
    .o(al_c4726cab));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_bdb3760b (
    .a(al_903070b1),
    .b(al_bfd664bf[0]),
    .c(al_bfd664bf[1]),
    .o(al_1308b999));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_971c58a1 (
    .a(al_69b84ba6[0]),
    .b(al_69b84ba6[1]),
    .c(al_69b84ba6[2]),
    .d(al_69b84ba6[3]),
    .e(al_69b84ba6[4]),
    .o(al_71fc1ad7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfffffffe7fffffff))
    al_51304b21 (
    .a(al_1308b999),
    .b(al_3014f961[0]),
    .c(al_3014f961[1]),
    .d(al_3014f961[2]),
    .e(al_3014f961[3]),
    .f(al_2ca0cac1),
    .o(al_8dcceed9));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1a403624 (
    .a(ddr_app_rdy),
    .b(al_cf00ed6f[4]),
    .c(al_5d3f410a[4]),
    .o(al_58fb4752[4]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_aaf28dc0 (
    .a(al_8dcceed9),
    .b(al_6db5b9d2),
    .c(al_3014f961[4]),
    .o(al_d1db9874[4]));
  AL_MAP_LUT5 #(
    .EQN("(~B*(D@(A*C*~(E)+~(A)*~(C)*E)))"),
    .INIT(32'h32011320))
    al_5b3caf58 (
    .a(al_1308b999),
    .b(al_6db5b9d2),
    .c(al_3014f961[0]),
    .d(al_3014f961[1]),
    .e(al_2ca0cac1),
    .o(al_d1db9874[1]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@C@A))"),
    .INIT(16'h2112))
    al_fe606af0 (
    .a(al_1308b999),
    .b(al_6db5b9d2),
    .c(al_3014f961[0]),
    .d(al_2ca0cac1),
    .o(al_d1db9874[0]));
  AL_MAP_LUT6 #(
    .EQN("(E@(~(A)*~(B)*~(C)*~(D)*~(F)+A*~(B)*~(C)*~(D)*~(F)+~(A)*B*~(C)*~(D)*~(F)+A*B*~(C)*~(D)*~(F)+~(A)*~(B)*C*~(D)*~(F)+A*~(B)*C*~(D)*~(F)+~(A)*B*C*~(D)*~(F)+A*B*C*~(D)*~(F)+~(A)*~(B)*~(C)*D*~(F)+A*~(B)*~(C)*D*~(F)+~(A)*B*~(C)*D*~(F)+A*B*~(C)*D*~(F)+~(A)*~(B)*C*D*~(F)+A*~(B)*C*D*~(F)+~(A)*B*C*D*~(F)+A*~(B)*~(C)*~(D)*F+~(A)*B*~(C)*~(D)*F+A*B*~(C)*~(D)*F+~(A)*~(B)*C*~(D)*F+A*~(B)*C*~(D)*F+~(A)*B*C*~(D)*F+A*B*C*~(D)*F+~(A)*~(B)*~(C)*D*F+A*~(B)*~(C)*D*F+~(A)*B*~(C)*D*F+A*B*~(C)*D*F+~(A)*~(B)*C*D*F+A*~(B)*C*D*F+~(A)*B*C*D*F+A*B*C*D*F))"),
    .INIT(64'h0001fffe80007fff))
    al_88ff0364 (
    .a(al_1308b999),
    .b(al_3014f961[0]),
    .c(al_3014f961[1]),
    .d(al_3014f961[2]),
    .e(al_3014f961[3]),
    .f(al_2ca0cac1),
    .o(al_adf8e398));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_4273b5ad (
    .a(al_adf8e398),
    .b(al_6db5b9d2),
    .o(al_d1db9874[3]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(E@(A*C*D*~(F)+~(A)*~(C)*~(D)*F)))"),
    .INIT(64'h3332000113332000))
    al_34c92c82 (
    .a(al_1308b999),
    .b(al_6db5b9d2),
    .c(al_3014f961[0]),
    .d(al_3014f961[1]),
    .e(al_3014f961[2]),
    .f(al_2ca0cac1),
    .o(al_d1db9874[2]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_3825ea48 (
    .a(al_d1db9874[4]),
    .b(al_d1db9874[3]),
    .c(al_d1db9874[1]),
    .d(al_d1db9874[0]),
    .e(al_d1db9874[2]),
    .o(al_355d4013));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(~C*A))"),
    .INIT(16'h39c6))
    al_1e40b4ed (
    .a(al_99c445b5[0]),
    .b(al_99c445b5[1]),
    .c(al_879aba03[0]),
    .d(al_879aba03[1]),
    .o(al_a9ec6721[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_7f17f864 (
    .a(al_2ee87d50),
    .b(al_b65fb56b),
    .c(al_40276cd4),
    .d(al_c4726cab),
    .o(al_e4f8f2fd));
  AL_MAP_LUT5 #(
    .EQN("(~E*~B*~A*~(D*C))"),
    .INIT(32'h00000111))
    al_973caf56 (
    .a(al_355d4013),
    .b(al_e4f8f2fd),
    .c(al_a7c937ec),
    .d(al_71fc1ad7),
    .e(al_69b84ba6[5]),
    .o(al_aab837cc));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_40143d1d (
    .a(al_903070b1),
    .b(al_bfd664bf[0]),
    .c(al_bfd664bf[1]),
    .o(al_a7c937ec));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*~B*~A)"),
    .INIT(32'h00000100))
    al_ccf88036 (
    .a(al_a9ec6721[1]),
    .b(al_58fb4752[3]),
    .c(al_58fb4752[4]),
    .d(init_calib_complete),
    .e(al_2d3f245b),
    .o(al_2ee87d50));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(~C*A))"),
    .INIT(16'h39c6))
    al_c5d7cba0 (
    .a(al_bd042336[0]),
    .b(al_bd042336[1]),
    .c(al_66e5f5b5[0]),
    .d(al_66e5f5b5[1]),
    .o(al_66006155));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*~A)"),
    .INIT(32'h00000400))
    al_a03f7360 (
    .a(al_66006155),
    .b(al_58fb4752[3]),
    .c(al_58fb4752[4]),
    .d(init_calib_complete),
    .e(al_7c9229ee),
    .o(al_b65fb56b));
  AL_DFF_0 al_8cad231 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aab837cc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rdy));
  AL_DFF_0 al_cd6c74c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[8]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[8]));
  AL_DFF_0 al_984a6f0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[9]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[9]));
  AL_DFF_0 al_a7d847fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[10]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[10]));
  AL_DFF_0 al_6a077416 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[11]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[11]));
  AL_DFF_0 al_d86303d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[12]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[12]));
  AL_DFF_0 al_ca9af6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[13]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[13]));
  AL_DFF_0 al_fe974a59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[14]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[14]));
  AL_DFF_0 al_f714a381 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[15]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[15]));
  AL_DFF_0 al_34fc6f60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[16]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[16]));
  AL_DFF_0 al_d0e760ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[17]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[17]));
  AL_DFF_0 al_45cdb76b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[18]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[18]));
  AL_DFF_0 al_8c96ade3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[19]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[19]));
  AL_DFF_0 al_f9714922 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[20]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[20]));
  AL_DFF_0 al_4ef1ef52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[21]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[21]));
  AL_DFF_0 al_6536e0f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[22]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[22]));
  AL_DFF_0 al_a7ee5a16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[23]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[23]));
  AL_DFF_0 al_5d1b5c9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[24]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[24]));
  AL_DFF_0 al_c26a6e44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[25]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[25]));
  AL_DFF_0 al_40f99812 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[26]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[26]));
  AL_DFF_0 al_9915760b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[3]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[3]));
  AL_DFF_0 al_70d938c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[4]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[4]));
  AL_DFF_0 al_11d6c91e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[5]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[5]));
  AL_DFF_0 al_27d204 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[6]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[6]));
  AL_DFF_0 al_2a27edcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_addr[7]),
    .en(al_e58efc01),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_cf00ed6f[7]));
  AL_DFF_0 al_f1238156 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[8]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[8]));
  AL_DFF_0 al_62e318ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[9]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[9]));
  AL_DFF_0 al_4bb89dcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[10]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[10]));
  AL_DFF_0 al_e02afadb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[11]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[11]));
  AL_DFF_0 al_182279b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[12]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[12]));
  AL_DFF_0 al_b2d9f5dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[13]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[13]));
  AL_DFF_0 al_723f1017 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[14]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[14]));
  AL_DFF_0 al_2eb1942c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[15]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[15]));
  AL_DFF_0 al_add88d57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[16]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[16]));
  AL_DFF_0 al_29f83867 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[17]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[17]));
  AL_DFF_0 al_bdd8eda6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[18]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[18]));
  AL_DFF_0 al_63c87a21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[19]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[19]));
  AL_DFF_0 al_b27662d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[20]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[20]));
  AL_DFF_0 al_5b215f8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[21]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[21]));
  AL_DFF_0 al_d3ba44c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[22]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[22]));
  AL_DFF_0 al_5087371b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[23]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[23]));
  AL_DFF_0 al_f22d206d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[24]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[24]));
  AL_DFF_0 al_a7782a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[25]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[25]));
  AL_DFF_0 al_ccd40957 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[26]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[26]));
  AL_DFF_0 al_e7e6da96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[3]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[3]));
  AL_DFF_0 al_56b82f21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[4]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[4]));
  AL_DFF_0 al_ce512569 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[5]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[5]));
  AL_DFF_0 al_487d8a3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[6]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[6]));
  AL_DFF_0 al_d89f5dc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf00ed6f[7]),
    .en(ddr_app_rdy),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5d3f410a[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_307e87a7 (
    .a(ddr_app_cmd[0]),
    .b(ddr_app_rdy),
    .c(al_65621cdc[0]),
    .o(al_7c29888a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_370a42ca (
    .a(ddr_app_cmd[1]),
    .b(ddr_app_rdy),
    .c(al_65621cdc[1]),
    .o(al_4c03fc24));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_511a1396 (
    .a(ddr_app_cmd[2]),
    .b(ddr_app_rdy),
    .c(al_65621cdc[2]),
    .o(al_330ee0e3));
  AL_DFF_0 al_3b1386df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c29888a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65621cdc[0]));
  AL_DFF_0 al_4f499322 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c03fc24),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65621cdc[1]));
  AL_DFF_0 al_de8222ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_330ee0e3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65621cdc[2]));
  AL_DFF_0 al_7b5aa2b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfd664bf[0]));
  AL_DFF_0 al_80e2a54b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfd664bf[1]));
  AL_DFF_0 al_cc1c67ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_88a8db2c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfd664bf[2]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_d43eacbd (
    .a(al_a56ffae1),
    .b(al_b2febcce[1]),
    .o(al_9c1746a1));
  AL_DFF_0 al_347edb75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9c1746a1),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(ddr_app_rd_data_end));
  AL_DFF_0 al_df43fcf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f33f7f41),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data_valid));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT(16'h1130))
    al_b7b7e02 (
    .a(al_f5b95ad4),
    .b(al_6db5b9d2),
    .c(ddr_app_rd_data_valid),
    .d(al_83931c3d),
    .o(al_f33f7f41));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_c9b1998 (
    .a(al_f5b95ad4),
    .b(al_70117344),
    .c(al_ebd79caa),
    .o(al_8c8985a1));
  AL_DFF_0 al_c3cce91f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c8985a1),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_3cc6b708));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_230efbfa (
    .i(al_3cc6b708),
    .o(al_13d66540));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_eeebd14 (
    .i(al_13d66540),
    .o(al_70117344));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_833abb0d (
    .i(al_4e8fb619),
    .o(al_da88ced7[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7390317a (
    .i(al_da88ced7[0]),
    .o(al_5b144427));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a086ba83 (
    .i(al_fd6a3ba4),
    .o(al_da88ced7[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a0af0316 (
    .i(al_da88ced7[1]),
    .o(al_42d963e6));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b0f2e981 (
    .i(al_b3cfcb5e),
    .o(al_da88ced7[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c330fe15 (
    .i(al_da88ced7[2]),
    .o(al_f1015bac));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c235c0f8 (
    .i(al_9a7b3b80),
    .o(al_da88ced7[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e31fd992 (
    .i(al_da88ced7[3]),
    .o(al_8cf002a4));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_6895256a (
    .a(al_880139ce[0]),
    .b(al_880139ce[1]),
    .c(al_880139ce[2]),
    .d(al_880139ce[3]),
    .e(al_880139ce[4]),
    .f(al_f1015bac),
    .o(al_adc73f46));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_8c11ba36 (
    .a(al_8e42692a[0]),
    .b(al_8e42692a[1]),
    .c(al_8e42692a[2]),
    .d(al_8e42692a[3]),
    .e(al_8e42692a[4]),
    .f(al_42d963e6),
    .o(al_2db7ae9f));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_58988e3d (
    .a(al_620ff4d8[0]),
    .b(al_620ff4d8[1]),
    .c(al_620ff4d8[2]),
    .d(al_620ff4d8[3]),
    .e(al_620ff4d8[4]),
    .f(al_5b144427),
    .o(al_4c1ffe8c));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_3205ba01 (
    .a(al_8119a127[0]),
    .b(al_8119a127[1]),
    .c(al_8119a127[2]),
    .d(al_8119a127[3]),
    .e(al_8119a127[4]),
    .f(al_8cf002a4),
    .o(al_99dca23));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_72e78a53 (
    .a(al_7905d584),
    .b(al_31a3e7af[192]),
    .c(al_955db046[192]),
    .o(al_f3aa16a9[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_57557980 (
    .a(al_7905d584),
    .b(al_31a3e7af[193]),
    .c(al_955db046[193]),
    .o(al_f3aa16a9[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f1eef774 (
    .a(al_7905d584),
    .b(al_31a3e7af[194]),
    .c(al_955db046[194]),
    .o(al_f3aa16a9[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9c3a3d37 (
    .a(al_7905d584),
    .b(al_31a3e7af[195]),
    .c(al_955db046[195]),
    .o(al_f3aa16a9[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ca47a7 (
    .a(al_7905d584),
    .b(al_31a3e7af[196]),
    .c(al_955db046[196]),
    .o(al_f3aa16a9[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5ad05f3d (
    .a(al_7905d584),
    .b(al_31a3e7af[197]),
    .c(al_955db046[197]),
    .o(al_f3aa16a9[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8a22bad9 (
    .a(al_ba6805c2),
    .b(al_31a3e7af[186]),
    .c(al_955db046[186]),
    .o(al_d0d403d6[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8849c9b (
    .a(al_ba6805c2),
    .b(al_31a3e7af[187]),
    .c(al_955db046[187]),
    .o(al_d0d403d6[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9e4b0191 (
    .a(al_ba6805c2),
    .b(al_31a3e7af[188]),
    .c(al_955db046[188]),
    .o(al_d0d403d6[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_77c1766a (
    .a(al_ba6805c2),
    .b(al_31a3e7af[189]),
    .c(al_955db046[189]),
    .o(al_d0d403d6[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ec4b5079 (
    .a(al_ba6805c2),
    .b(al_31a3e7af[190]),
    .c(al_955db046[190]),
    .o(al_d0d403d6[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_32baac27 (
    .a(al_ba6805c2),
    .b(al_31a3e7af[191]),
    .c(al_955db046[191]),
    .o(al_d0d403d6[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b3211e67 (
    .a(al_957b61e0),
    .b(al_31a3e7af[180]),
    .c(al_955db046[180]),
    .o(al_2c2ca002[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fb0c8540 (
    .a(al_957b61e0),
    .b(al_31a3e7af[181]),
    .c(al_955db046[181]),
    .o(al_2c2ca002[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d385467a (
    .a(al_957b61e0),
    .b(al_31a3e7af[182]),
    .c(al_955db046[182]),
    .o(al_2c2ca002[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ccf2c355 (
    .a(al_957b61e0),
    .b(al_31a3e7af[183]),
    .c(al_955db046[183]),
    .o(al_2c2ca002[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_606d94f7 (
    .a(al_957b61e0),
    .b(al_31a3e7af[184]),
    .c(al_955db046[184]),
    .o(al_2c2ca002[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b2b20fa6 (
    .a(al_957b61e0),
    .b(al_31a3e7af[185]),
    .c(al_955db046[185]),
    .o(al_2c2ca002[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2dbcf81b (
    .a(al_9e2fe654),
    .b(al_31a3e7af[174]),
    .c(al_955db046[174]),
    .o(al_5c25a985[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_faf1a489 (
    .a(al_9e2fe654),
    .b(al_31a3e7af[175]),
    .c(al_955db046[175]),
    .o(al_5c25a985[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3aa4dc3d (
    .a(al_9e2fe654),
    .b(al_31a3e7af[176]),
    .c(al_955db046[176]),
    .o(al_5c25a985[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a724a21d (
    .a(al_9e2fe654),
    .b(al_31a3e7af[177]),
    .c(al_955db046[177]),
    .o(al_5c25a985[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_10cc59bd (
    .a(al_9e2fe654),
    .b(al_31a3e7af[178]),
    .c(al_955db046[178]),
    .o(al_5c25a985[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e22e573e (
    .a(al_9e2fe654),
    .b(al_31a3e7af[179]),
    .c(al_955db046[179]),
    .o(al_5c25a985[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f5d4ff09 (
    .a(al_2cac5213),
    .b(al_31a3e7af[168]),
    .c(al_955db046[168]),
    .o(al_8b88a45c[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_73091e85 (
    .a(al_2cac5213),
    .b(al_31a3e7af[169]),
    .c(al_955db046[169]),
    .o(al_8b88a45c[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9c8fe9d9 (
    .a(al_2cac5213),
    .b(al_31a3e7af[170]),
    .c(al_955db046[170]),
    .o(al_8b88a45c[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_20a8a465 (
    .a(al_2cac5213),
    .b(al_31a3e7af[171]),
    .c(al_955db046[171]),
    .o(al_8b88a45c[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c14deebf (
    .a(al_2cac5213),
    .b(al_31a3e7af[172]),
    .c(al_955db046[172]),
    .o(al_8b88a45c[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7b3b4bdc (
    .a(al_2cac5213),
    .b(al_31a3e7af[173]),
    .c(al_955db046[173]),
    .o(al_8b88a45c[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a1e4c1f8 (
    .a(al_c5c99a19),
    .b(al_31a3e7af[162]),
    .c(al_955db046[162]),
    .o(al_d88fcc0f[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_68237ce (
    .a(al_c5c99a19),
    .b(al_31a3e7af[163]),
    .c(al_955db046[163]),
    .o(al_d88fcc0f[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_12ae5ff5 (
    .a(al_c5c99a19),
    .b(al_31a3e7af[164]),
    .c(al_955db046[164]),
    .o(al_d88fcc0f[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6bbdfeef (
    .a(al_c5c99a19),
    .b(al_31a3e7af[165]),
    .c(al_955db046[165]),
    .o(al_d88fcc0f[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ca50d0df (
    .a(al_c5c99a19),
    .b(al_31a3e7af[166]),
    .c(al_955db046[166]),
    .o(al_d88fcc0f[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f5602d40 (
    .a(al_c5c99a19),
    .b(al_31a3e7af[167]),
    .c(al_955db046[167]),
    .o(al_d88fcc0f[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_28cff8ab (
    .a(al_9b71a4e4),
    .b(al_31a3e7af[156]),
    .c(al_955db046[156]),
    .o(al_b8da42f7[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2a06cb70 (
    .a(al_9b71a4e4),
    .b(al_31a3e7af[157]),
    .c(al_955db046[157]),
    .o(al_b8da42f7[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f1a9d2f2 (
    .a(al_9b71a4e4),
    .b(al_31a3e7af[158]),
    .c(al_955db046[158]),
    .o(al_b8da42f7[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4518573e (
    .a(al_9b71a4e4),
    .b(al_31a3e7af[159]),
    .c(al_955db046[159]),
    .o(al_b8da42f7[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_40da0370 (
    .a(al_9b71a4e4),
    .b(al_31a3e7af[160]),
    .c(al_955db046[160]),
    .o(al_b8da42f7[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_212dd592 (
    .a(al_9b71a4e4),
    .b(al_31a3e7af[161]),
    .c(al_955db046[161]),
    .o(al_b8da42f7[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8b2890ee (
    .a(al_312b2dca),
    .b(al_31a3e7af[150]),
    .c(al_955db046[150]),
    .o(al_f033fc44[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_95c6db9b (
    .a(al_312b2dca),
    .b(al_31a3e7af[151]),
    .c(al_955db046[151]),
    .o(al_f033fc44[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_386464e1 (
    .a(al_312b2dca),
    .b(al_31a3e7af[152]),
    .c(al_955db046[152]),
    .o(al_f033fc44[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_56cc95c5 (
    .a(al_312b2dca),
    .b(al_31a3e7af[153]),
    .c(al_955db046[153]),
    .o(al_f033fc44[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b844667c (
    .a(al_312b2dca),
    .b(al_31a3e7af[154]),
    .c(al_955db046[154]),
    .o(al_f033fc44[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_71472b2d (
    .a(al_312b2dca),
    .b(al_31a3e7af[155]),
    .c(al_955db046[155]),
    .o(al_f033fc44[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bfee1ad1 (
    .a(al_b49bcb3),
    .b(al_31a3e7af[144]),
    .c(al_955db046[144]),
    .o(al_3a9b666[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ced01884 (
    .a(al_b49bcb3),
    .b(al_31a3e7af[145]),
    .c(al_955db046[145]),
    .o(al_3a9b666[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ddc033d8 (
    .a(al_b49bcb3),
    .b(al_31a3e7af[146]),
    .c(al_955db046[146]),
    .o(al_3a9b666[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_58c7f678 (
    .a(al_b49bcb3),
    .b(al_31a3e7af[147]),
    .c(al_955db046[147]),
    .o(al_3a9b666[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_cd27e42e (
    .a(al_b49bcb3),
    .b(al_31a3e7af[148]),
    .c(al_955db046[148]),
    .o(al_3a9b666[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_553c5d9d (
    .a(al_b49bcb3),
    .b(al_31a3e7af[149]),
    .c(al_955db046[149]),
    .o(al_3a9b666[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2424ba0a (
    .a(al_d8d52ddc),
    .b(al_31a3e7af[138]),
    .c(al_955db046[138]),
    .o(al_a5ad4b3c[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_79b8623d (
    .a(al_d8d52ddc),
    .b(al_31a3e7af[139]),
    .c(al_955db046[139]),
    .o(al_a5ad4b3c[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5ebd4720 (
    .a(al_d8d52ddc),
    .b(al_31a3e7af[140]),
    .c(al_955db046[140]),
    .o(al_a5ad4b3c[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b9aa3e27 (
    .a(al_d8d52ddc),
    .b(al_31a3e7af[141]),
    .c(al_955db046[141]),
    .o(al_a5ad4b3c[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5ae2462b (
    .a(al_d8d52ddc),
    .b(al_31a3e7af[142]),
    .c(al_955db046[142]),
    .o(al_a5ad4b3c[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_54f54613 (
    .a(al_d8d52ddc),
    .b(al_31a3e7af[143]),
    .c(al_955db046[143]),
    .o(al_a5ad4b3c[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c4b4a580 (
    .a(al_3ed1abca),
    .b(al_31a3e7af[246]),
    .c(al_955db046[246]),
    .o(al_a3fa002d[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_cde12767 (
    .a(al_3ed1abca),
    .b(al_31a3e7af[247]),
    .c(al_955db046[247]),
    .o(al_a3fa002d[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8e4d7e1e (
    .a(al_3ed1abca),
    .b(al_31a3e7af[248]),
    .c(al_955db046[248]),
    .o(al_a3fa002d[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b0a72ba (
    .a(al_3ed1abca),
    .b(al_31a3e7af[249]),
    .c(al_955db046[249]),
    .o(al_a3fa002d[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6c724d33 (
    .a(al_3ed1abca),
    .b(al_31a3e7af[250]),
    .c(al_955db046[250]),
    .o(al_a3fa002d[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_43cd2a91 (
    .a(al_3ed1abca),
    .b(al_31a3e7af[251]),
    .c(al_955db046[251]),
    .o(al_a3fa002d[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ab70f99f (
    .a(al_f07cc0e),
    .b(al_31a3e7af[132]),
    .c(al_955db046[132]),
    .o(al_b9ca6681[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8515e66e (
    .a(al_f07cc0e),
    .b(al_31a3e7af[133]),
    .c(al_955db046[133]),
    .o(al_b9ca6681[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ff745029 (
    .a(al_f07cc0e),
    .b(al_31a3e7af[134]),
    .c(al_955db046[134]),
    .o(al_b9ca6681[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ef706d25 (
    .a(al_f07cc0e),
    .b(al_31a3e7af[135]),
    .c(al_955db046[135]),
    .o(al_b9ca6681[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c78d1f05 (
    .a(al_f07cc0e),
    .b(al_31a3e7af[136]),
    .c(al_955db046[136]),
    .o(al_b9ca6681[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_cd000fea (
    .a(al_f07cc0e),
    .b(al_31a3e7af[137]),
    .c(al_955db046[137]),
    .o(al_b9ca6681[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bd4beee3 (
    .a(al_a4c76fab),
    .b(al_31a3e7af[126]),
    .c(al_955db046[126]),
    .o(al_69204309[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5daf4807 (
    .a(al_a4c76fab),
    .b(al_31a3e7af[127]),
    .c(al_955db046[127]),
    .o(al_69204309[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_eaa45b6c (
    .a(al_a4c76fab),
    .b(al_31a3e7af[128]),
    .c(al_955db046[128]),
    .o(al_69204309[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c66efa94 (
    .a(al_a4c76fab),
    .b(al_31a3e7af[129]),
    .c(al_955db046[129]),
    .o(al_69204309[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_713d089f (
    .a(al_a4c76fab),
    .b(al_31a3e7af[130]),
    .c(al_955db046[130]),
    .o(al_69204309[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5c52017d (
    .a(al_a4c76fab),
    .b(al_31a3e7af[131]),
    .c(al_955db046[131]),
    .o(al_69204309[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1e8f89b3 (
    .a(al_ad24301),
    .b(al_31a3e7af[120]),
    .c(al_955db046[120]),
    .o(al_98058573[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_af4c949a (
    .a(al_ad24301),
    .b(al_31a3e7af[121]),
    .c(al_955db046[121]),
    .o(al_98058573[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e83a7085 (
    .a(al_ad24301),
    .b(al_31a3e7af[122]),
    .c(al_955db046[122]),
    .o(al_98058573[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8936f9c8 (
    .a(al_ad24301),
    .b(al_31a3e7af[123]),
    .c(al_955db046[123]),
    .o(al_98058573[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5c2b2656 (
    .a(al_ad24301),
    .b(al_31a3e7af[124]),
    .c(al_955db046[124]),
    .o(al_98058573[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b0a83f2c (
    .a(al_ad24301),
    .b(al_31a3e7af[125]),
    .c(al_955db046[125]),
    .o(al_98058573[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_55c2fd7d (
    .a(al_8091f068),
    .b(al_31a3e7af[114]),
    .c(al_955db046[114]),
    .o(al_63020263[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e7154d56 (
    .a(al_8091f068),
    .b(al_31a3e7af[115]),
    .c(al_955db046[115]),
    .o(al_63020263[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4707c86f (
    .a(al_8091f068),
    .b(al_31a3e7af[116]),
    .c(al_955db046[116]),
    .o(al_63020263[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6b9fb489 (
    .a(al_8091f068),
    .b(al_31a3e7af[117]),
    .c(al_955db046[117]),
    .o(al_63020263[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2d9af3b4 (
    .a(al_8091f068),
    .b(al_31a3e7af[118]),
    .c(al_955db046[118]),
    .o(al_63020263[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d6092f2f (
    .a(al_8091f068),
    .b(al_31a3e7af[119]),
    .c(al_955db046[119]),
    .o(al_63020263[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3388895c (
    .a(al_af74714f),
    .b(al_31a3e7af[108]),
    .c(al_955db046[108]),
    .o(al_b7a189[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_491933d7 (
    .a(al_af74714f),
    .b(al_31a3e7af[109]),
    .c(al_955db046[109]),
    .o(al_b7a189[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f8936482 (
    .a(al_af74714f),
    .b(al_31a3e7af[110]),
    .c(al_955db046[110]),
    .o(al_b7a189[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b6487a4e (
    .a(al_af74714f),
    .b(al_31a3e7af[111]),
    .c(al_955db046[111]),
    .o(al_b7a189[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f86f39f1 (
    .a(al_af74714f),
    .b(al_31a3e7af[112]),
    .c(al_955db046[112]),
    .o(al_b7a189[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d3f0ed5f (
    .a(al_af74714f),
    .b(al_31a3e7af[113]),
    .c(al_955db046[113]),
    .o(al_b7a189[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2488b76c (
    .a(al_3310bf9b),
    .b(al_31a3e7af[102]),
    .c(al_955db046[102]),
    .o(al_c527aa4e[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b28afd99 (
    .a(al_3310bf9b),
    .b(al_31a3e7af[103]),
    .c(al_955db046[103]),
    .o(al_c527aa4e[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7e0c8d00 (
    .a(al_3310bf9b),
    .b(al_31a3e7af[104]),
    .c(al_955db046[104]),
    .o(al_c527aa4e[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9c497581 (
    .a(al_3310bf9b),
    .b(al_31a3e7af[105]),
    .c(al_955db046[105]),
    .o(al_c527aa4e[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_58917b28 (
    .a(al_3310bf9b),
    .b(al_31a3e7af[106]),
    .c(al_955db046[106]),
    .o(al_c527aa4e[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_34d82824 (
    .a(al_3310bf9b),
    .b(al_31a3e7af[107]),
    .c(al_955db046[107]),
    .o(al_c527aa4e[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_23270d18 (
    .a(al_a6167193),
    .b(al_31a3e7af[96]),
    .c(al_955db046[96]),
    .o(al_407652d9[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4df4d3b3 (
    .a(al_a6167193),
    .b(al_31a3e7af[97]),
    .c(al_955db046[97]),
    .o(al_407652d9[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_843f538 (
    .a(al_a6167193),
    .b(al_31a3e7af[98]),
    .c(al_955db046[98]),
    .o(al_407652d9[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b14fc8d0 (
    .a(al_a6167193),
    .b(al_31a3e7af[99]),
    .c(al_955db046[99]),
    .o(al_407652d9[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8114c22a (
    .a(al_a6167193),
    .b(al_31a3e7af[100]),
    .c(al_955db046[100]),
    .o(al_407652d9[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e5d533c (
    .a(al_a6167193),
    .b(al_31a3e7af[101]),
    .c(al_955db046[101]),
    .o(al_407652d9[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_894ab772 (
    .a(al_3728ce00),
    .b(al_31a3e7af[90]),
    .c(al_955db046[90]),
    .o(al_fce7b5a9[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_16ec9a3a (
    .a(al_3728ce00),
    .b(al_31a3e7af[91]),
    .c(al_955db046[91]),
    .o(al_fce7b5a9[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3f9c61c4 (
    .a(al_3728ce00),
    .b(al_31a3e7af[92]),
    .c(al_955db046[92]),
    .o(al_fce7b5a9[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6be285de (
    .a(al_3728ce00),
    .b(al_31a3e7af[93]),
    .c(al_955db046[93]),
    .o(al_fce7b5a9[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6ede44e6 (
    .a(al_3728ce00),
    .b(al_31a3e7af[94]),
    .c(al_955db046[94]),
    .o(al_fce7b5a9[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ce8b014e (
    .a(al_3728ce00),
    .b(al_31a3e7af[95]),
    .c(al_955db046[95]),
    .o(al_fce7b5a9[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b8f8bbdc (
    .a(al_fd1400b6),
    .b(al_31a3e7af[84]),
    .c(al_955db046[84]),
    .o(al_87305132[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2b51ecce (
    .a(al_fd1400b6),
    .b(al_31a3e7af[85]),
    .c(al_955db046[85]),
    .o(al_87305132[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4076402d (
    .a(al_fd1400b6),
    .b(al_31a3e7af[86]),
    .c(al_955db046[86]),
    .o(al_87305132[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fd9af723 (
    .a(al_fd1400b6),
    .b(al_31a3e7af[87]),
    .c(al_955db046[87]),
    .o(al_87305132[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3a01669b (
    .a(al_fd1400b6),
    .b(al_31a3e7af[88]),
    .c(al_955db046[88]),
    .o(al_87305132[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1c49e452 (
    .a(al_fd1400b6),
    .b(al_31a3e7af[89]),
    .c(al_955db046[89]),
    .o(al_87305132[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_49554910 (
    .a(al_72450658),
    .b(al_31a3e7af[78]),
    .c(al_955db046[78]),
    .o(al_ed19afe1[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_471969f2 (
    .a(al_72450658),
    .b(al_31a3e7af[79]),
    .c(al_955db046[79]),
    .o(al_ed19afe1[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9e1c43f9 (
    .a(al_72450658),
    .b(al_31a3e7af[80]),
    .c(al_955db046[80]),
    .o(al_ed19afe1[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fbeb9269 (
    .a(al_72450658),
    .b(al_31a3e7af[81]),
    .c(al_955db046[81]),
    .o(al_ed19afe1[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e9a8a900 (
    .a(al_72450658),
    .b(al_31a3e7af[82]),
    .c(al_955db046[82]),
    .o(al_ed19afe1[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f3f89d57 (
    .a(al_72450658),
    .b(al_31a3e7af[83]),
    .c(al_955db046[83]),
    .o(al_ed19afe1[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_64884b9d (
    .a(al_733e11d7),
    .b(al_31a3e7af[240]),
    .c(al_955db046[240]),
    .o(al_77d19440[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bce82d16 (
    .a(al_733e11d7),
    .b(al_31a3e7af[241]),
    .c(al_955db046[241]),
    .o(al_77d19440[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bbc44a0 (
    .a(al_733e11d7),
    .b(al_31a3e7af[242]),
    .c(al_955db046[242]),
    .o(al_77d19440[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e1e5323a (
    .a(al_733e11d7),
    .b(al_31a3e7af[243]),
    .c(al_955db046[243]),
    .o(al_77d19440[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5b30ee59 (
    .a(al_733e11d7),
    .b(al_31a3e7af[244]),
    .c(al_955db046[244]),
    .o(al_77d19440[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ebf1dadd (
    .a(al_733e11d7),
    .b(al_31a3e7af[245]),
    .c(al_955db046[245]),
    .o(al_77d19440[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e5e9a9bd (
    .a(al_2c66a236),
    .b(al_31a3e7af[72]),
    .c(al_955db046[72]),
    .o(al_33614149[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2817b987 (
    .a(al_2c66a236),
    .b(al_31a3e7af[73]),
    .c(al_955db046[73]),
    .o(al_33614149[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d4e78c54 (
    .a(al_2c66a236),
    .b(al_31a3e7af[74]),
    .c(al_955db046[74]),
    .o(al_33614149[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_65f29f89 (
    .a(al_2c66a236),
    .b(al_31a3e7af[75]),
    .c(al_955db046[75]),
    .o(al_33614149[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_48be37dc (
    .a(al_2c66a236),
    .b(al_31a3e7af[76]),
    .c(al_955db046[76]),
    .o(al_33614149[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_db802c3a (
    .a(al_2c66a236),
    .b(al_31a3e7af[77]),
    .c(al_955db046[77]),
    .o(al_33614149[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c9343bf3 (
    .a(al_e3e65c55),
    .b(al_31a3e7af[66]),
    .c(al_955db046[66]),
    .o(al_175c7e02[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f3924437 (
    .a(al_e3e65c55),
    .b(al_31a3e7af[67]),
    .c(al_955db046[67]),
    .o(al_175c7e02[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_17bd7ee3 (
    .a(al_e3e65c55),
    .b(al_31a3e7af[68]),
    .c(al_955db046[68]),
    .o(al_175c7e02[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b504e5ce (
    .a(al_e3e65c55),
    .b(al_31a3e7af[69]),
    .c(al_955db046[69]),
    .o(al_175c7e02[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a6f5a673 (
    .a(al_e3e65c55),
    .b(al_31a3e7af[70]),
    .c(al_955db046[70]),
    .o(al_175c7e02[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d0a8c5fa (
    .a(al_e3e65c55),
    .b(al_31a3e7af[71]),
    .c(al_955db046[71]),
    .o(al_175c7e02[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_85a10f0 (
    .a(al_2eb834f5),
    .b(al_31a3e7af[60]),
    .c(al_955db046[60]),
    .o(al_b48e0e9a[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5f0454d4 (
    .a(al_2eb834f5),
    .b(al_31a3e7af[61]),
    .c(al_955db046[61]),
    .o(al_b48e0e9a[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8ab15172 (
    .a(al_2eb834f5),
    .b(al_31a3e7af[62]),
    .c(al_955db046[62]),
    .o(al_b48e0e9a[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3b7a70fc (
    .a(al_2eb834f5),
    .b(al_31a3e7af[63]),
    .c(al_955db046[63]),
    .o(al_b48e0e9a[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_42db083c (
    .a(al_2eb834f5),
    .b(al_31a3e7af[64]),
    .c(al_955db046[64]),
    .o(al_b48e0e9a[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_125b0199 (
    .a(al_2eb834f5),
    .b(al_31a3e7af[65]),
    .c(al_955db046[65]),
    .o(al_b48e0e9a[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2316721e (
    .a(al_ec10e78f),
    .b(al_31a3e7af[54]),
    .c(al_955db046[54]),
    .o(al_92e7eeea[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_caa7a613 (
    .a(al_ec10e78f),
    .b(al_31a3e7af[55]),
    .c(al_955db046[55]),
    .o(al_92e7eeea[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_436ca5b1 (
    .a(al_ec10e78f),
    .b(al_31a3e7af[56]),
    .c(al_955db046[56]),
    .o(al_92e7eeea[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_dc349e09 (
    .a(al_ec10e78f),
    .b(al_31a3e7af[57]),
    .c(al_955db046[57]),
    .o(al_92e7eeea[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2301d60a (
    .a(al_ec10e78f),
    .b(al_31a3e7af[58]),
    .c(al_955db046[58]),
    .o(al_92e7eeea[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_61183780 (
    .a(al_ec10e78f),
    .b(al_31a3e7af[59]),
    .c(al_955db046[59]),
    .o(al_92e7eeea[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e18523f3 (
    .a(al_e75d67c1),
    .b(al_31a3e7af[48]),
    .c(al_955db046[48]),
    .o(al_a6a612a6[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_598071e4 (
    .a(al_e75d67c1),
    .b(al_31a3e7af[49]),
    .c(al_955db046[49]),
    .o(al_a6a612a6[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b25681e7 (
    .a(al_e75d67c1),
    .b(al_31a3e7af[50]),
    .c(al_955db046[50]),
    .o(al_a6a612a6[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5b809d34 (
    .a(al_e75d67c1),
    .b(al_31a3e7af[51]),
    .c(al_955db046[51]),
    .o(al_a6a612a6[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_94649496 (
    .a(al_e75d67c1),
    .b(al_31a3e7af[52]),
    .c(al_955db046[52]),
    .o(al_a6a612a6[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d7f387ae (
    .a(al_e75d67c1),
    .b(al_31a3e7af[53]),
    .c(al_955db046[53]),
    .o(al_a6a612a6[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d176c0d8 (
    .a(al_316d230a),
    .b(al_31a3e7af[42]),
    .c(al_955db046[42]),
    .o(al_9427b946[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1bb297a5 (
    .a(al_316d230a),
    .b(al_31a3e7af[43]),
    .c(al_955db046[43]),
    .o(al_9427b946[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4e30293f (
    .a(al_316d230a),
    .b(al_31a3e7af[44]),
    .c(al_955db046[44]),
    .o(al_9427b946[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ba790e40 (
    .a(al_316d230a),
    .b(al_31a3e7af[45]),
    .c(al_955db046[45]),
    .o(al_9427b946[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c125110e (
    .a(al_316d230a),
    .b(al_31a3e7af[46]),
    .c(al_955db046[46]),
    .o(al_9427b946[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_38e58735 (
    .a(al_316d230a),
    .b(al_31a3e7af[47]),
    .c(al_955db046[47]),
    .o(al_9427b946[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b0c1f598 (
    .a(al_6d6f3341),
    .b(al_31a3e7af[36]),
    .c(al_955db046[36]),
    .o(al_9bc4f0be[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_80cb5fac (
    .a(al_6d6f3341),
    .b(al_31a3e7af[37]),
    .c(al_955db046[37]),
    .o(al_9bc4f0be[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_10fb09dc (
    .a(al_6d6f3341),
    .b(al_31a3e7af[38]),
    .c(al_955db046[38]),
    .o(al_9bc4f0be[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_34795402 (
    .a(al_6d6f3341),
    .b(al_31a3e7af[39]),
    .c(al_955db046[39]),
    .o(al_9bc4f0be[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b2cfcca2 (
    .a(al_6d6f3341),
    .b(al_31a3e7af[40]),
    .c(al_955db046[40]),
    .o(al_9bc4f0be[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b18f2fa0 (
    .a(al_6d6f3341),
    .b(al_31a3e7af[41]),
    .c(al_955db046[41]),
    .o(al_9bc4f0be[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_777e72fd (
    .a(al_898acbc2),
    .b(al_31a3e7af[30]),
    .c(al_955db046[30]),
    .o(al_764d3602[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8432c85b (
    .a(al_898acbc2),
    .b(al_31a3e7af[31]),
    .c(al_955db046[31]),
    .o(al_764d3602[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_36cd0c00 (
    .a(al_898acbc2),
    .b(al_31a3e7af[32]),
    .c(al_955db046[32]),
    .o(al_764d3602[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_91a89c9a (
    .a(al_898acbc2),
    .b(al_31a3e7af[33]),
    .c(al_955db046[33]),
    .o(al_764d3602[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b063adb2 (
    .a(al_898acbc2),
    .b(al_31a3e7af[34]),
    .c(al_955db046[34]),
    .o(al_764d3602[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3ec6c882 (
    .a(al_898acbc2),
    .b(al_31a3e7af[35]),
    .c(al_955db046[35]),
    .o(al_764d3602[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_74733827 (
    .a(al_e1d70a3d),
    .b(al_31a3e7af[24]),
    .c(al_955db046[24]),
    .o(al_5a84549[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_86feec30 (
    .a(al_e1d70a3d),
    .b(al_31a3e7af[25]),
    .c(al_955db046[25]),
    .o(al_5a84549[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e05c1aa (
    .a(al_e1d70a3d),
    .b(al_31a3e7af[26]),
    .c(al_955db046[26]),
    .o(al_5a84549[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ab568f70 (
    .a(al_e1d70a3d),
    .b(al_31a3e7af[27]),
    .c(al_955db046[27]),
    .o(al_5a84549[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d463679e (
    .a(al_e1d70a3d),
    .b(al_31a3e7af[28]),
    .c(al_955db046[28]),
    .o(al_5a84549[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_507bbafc (
    .a(al_e1d70a3d),
    .b(al_31a3e7af[29]),
    .c(al_955db046[29]),
    .o(al_5a84549[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2ef49c47 (
    .a(al_fdf8d449),
    .b(al_31a3e7af[18]),
    .c(al_955db046[18]),
    .o(al_e5342096[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e82db760 (
    .a(al_fdf8d449),
    .b(al_31a3e7af[19]),
    .c(al_955db046[19]),
    .o(al_e5342096[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b6ecdd5 (
    .a(al_fdf8d449),
    .b(al_31a3e7af[20]),
    .c(al_955db046[20]),
    .o(al_e5342096[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8c593201 (
    .a(al_fdf8d449),
    .b(al_31a3e7af[21]),
    .c(al_955db046[21]),
    .o(al_e5342096[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7abfc787 (
    .a(al_fdf8d449),
    .b(al_31a3e7af[22]),
    .c(al_955db046[22]),
    .o(al_e5342096[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_45aad212 (
    .a(al_fdf8d449),
    .b(al_31a3e7af[23]),
    .c(al_955db046[23]),
    .o(al_e5342096[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_cfd593a2 (
    .a(al_6aad2723),
    .b(al_31a3e7af[234]),
    .c(al_955db046[234]),
    .o(al_98c6a23b[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_de41d659 (
    .a(al_6aad2723),
    .b(al_31a3e7af[235]),
    .c(al_955db046[235]),
    .o(al_98c6a23b[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_423d9f8d (
    .a(al_6aad2723),
    .b(al_31a3e7af[236]),
    .c(al_955db046[236]),
    .o(al_98c6a23b[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_706dc6ef (
    .a(al_6aad2723),
    .b(al_31a3e7af[237]),
    .c(al_955db046[237]),
    .o(al_98c6a23b[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_89e83e2c (
    .a(al_6aad2723),
    .b(al_31a3e7af[238]),
    .c(al_955db046[238]),
    .o(al_98c6a23b[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_81f22266 (
    .a(al_6aad2723),
    .b(al_31a3e7af[239]),
    .c(al_955db046[239]),
    .o(al_98c6a23b[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_aead4397 (
    .a(al_be012e15),
    .b(al_31a3e7af[12]),
    .c(al_955db046[12]),
    .o(al_27ec7185[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a63a91b4 (
    .a(al_be012e15),
    .b(al_31a3e7af[13]),
    .c(al_955db046[13]),
    .o(al_27ec7185[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4e347a49 (
    .a(al_be012e15),
    .b(al_31a3e7af[14]),
    .c(al_955db046[14]),
    .o(al_27ec7185[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2004d80 (
    .a(al_be012e15),
    .b(al_31a3e7af[15]),
    .c(al_955db046[15]),
    .o(al_27ec7185[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3111f793 (
    .a(al_be012e15),
    .b(al_31a3e7af[16]),
    .c(al_955db046[16]),
    .o(al_27ec7185[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ae9ec90a (
    .a(al_be012e15),
    .b(al_31a3e7af[17]),
    .c(al_955db046[17]),
    .o(al_27ec7185[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f23f22ba (
    .a(al_3bfb38e8),
    .b(al_31a3e7af[6]),
    .c(al_955db046[6]),
    .o(al_ea67686c[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_73e28ad5 (
    .a(al_3bfb38e8),
    .b(al_31a3e7af[7]),
    .c(al_955db046[7]),
    .o(al_ea67686c[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4d2f670c (
    .a(al_3bfb38e8),
    .b(al_31a3e7af[8]),
    .c(al_955db046[8]),
    .o(al_ea67686c[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d8d6e06 (
    .a(al_3bfb38e8),
    .b(al_31a3e7af[9]),
    .c(al_955db046[9]),
    .o(al_ea67686c[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fb5ed9f (
    .a(al_3bfb38e8),
    .b(al_31a3e7af[10]),
    .c(al_955db046[10]),
    .o(al_ea67686c[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d0681a75 (
    .a(al_3bfb38e8),
    .b(al_31a3e7af[11]),
    .c(al_955db046[11]),
    .o(al_ea67686c[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5fec3d91 (
    .a(al_d2cdc7c9),
    .b(al_31a3e7af[0]),
    .c(al_955db046[0]),
    .o(al_b04b1b3b[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a5267053 (
    .a(al_d2cdc7c9),
    .b(al_31a3e7af[1]),
    .c(al_955db046[1]),
    .o(al_b04b1b3b[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_69e795e1 (
    .a(al_d2cdc7c9),
    .b(al_31a3e7af[2]),
    .c(al_955db046[2]),
    .o(al_b04b1b3b[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_686be75d (
    .a(al_d2cdc7c9),
    .b(al_31a3e7af[3]),
    .c(al_955db046[3]),
    .o(al_b04b1b3b[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e5b17e4b (
    .a(al_d2cdc7c9),
    .b(al_31a3e7af[4]),
    .c(al_955db046[4]),
    .o(al_b04b1b3b[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1d81af4a (
    .a(al_d2cdc7c9),
    .b(al_31a3e7af[5]),
    .c(al_955db046[5]),
    .o(al_b04b1b3b[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7bc57faf (
    .a(al_84ac14c0),
    .b(al_31a3e7af[228]),
    .c(al_955db046[228]),
    .o(al_c0d076bb[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ec7913cd (
    .a(al_84ac14c0),
    .b(al_31a3e7af[229]),
    .c(al_955db046[229]),
    .o(al_c0d076bb[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2d282da7 (
    .a(al_84ac14c0),
    .b(al_31a3e7af[230]),
    .c(al_955db046[230]),
    .o(al_c0d076bb[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3ab79fbb (
    .a(al_84ac14c0),
    .b(al_31a3e7af[231]),
    .c(al_955db046[231]),
    .o(al_c0d076bb[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f9fb2ce1 (
    .a(al_84ac14c0),
    .b(al_31a3e7af[232]),
    .c(al_955db046[232]),
    .o(al_c0d076bb[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2138c7ad (
    .a(al_84ac14c0),
    .b(al_31a3e7af[233]),
    .c(al_955db046[233]),
    .o(al_c0d076bb[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3ed8680c (
    .a(al_1b504c84),
    .b(al_31a3e7af[222]),
    .c(al_955db046[222]),
    .o(al_d55b2543[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_56f8e2c2 (
    .a(al_1b504c84),
    .b(al_31a3e7af[223]),
    .c(al_955db046[223]),
    .o(al_d55b2543[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a2642a02 (
    .a(al_1b504c84),
    .b(al_31a3e7af[224]),
    .c(al_955db046[224]),
    .o(al_d55b2543[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f16bd1d3 (
    .a(al_1b504c84),
    .b(al_31a3e7af[225]),
    .c(al_955db046[225]),
    .o(al_d55b2543[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b58df164 (
    .a(al_1b504c84),
    .b(al_31a3e7af[226]),
    .c(al_955db046[226]),
    .o(al_d55b2543[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5d2aa827 (
    .a(al_1b504c84),
    .b(al_31a3e7af[227]),
    .c(al_955db046[227]),
    .o(al_d55b2543[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c3041bce (
    .a(al_a6be8738),
    .b(al_31a3e7af[216]),
    .c(al_955db046[216]),
    .o(al_5577a41[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_24840f54 (
    .a(al_a6be8738),
    .b(al_31a3e7af[217]),
    .c(al_955db046[217]),
    .o(al_5577a41[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_605a7bad (
    .a(al_a6be8738),
    .b(al_31a3e7af[218]),
    .c(al_955db046[218]),
    .o(al_5577a41[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_909fe858 (
    .a(al_a6be8738),
    .b(al_31a3e7af[219]),
    .c(al_955db046[219]),
    .o(al_5577a41[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c412b012 (
    .a(al_a6be8738),
    .b(al_31a3e7af[220]),
    .c(al_955db046[220]),
    .o(al_5577a41[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c3685ef (
    .a(al_a6be8738),
    .b(al_31a3e7af[221]),
    .c(al_955db046[221]),
    .o(al_5577a41[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_81cadeb8 (
    .a(al_c21b49ee),
    .b(al_31a3e7af[210]),
    .c(al_955db046[210]),
    .o(al_b0408eb[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2c8d6b00 (
    .a(al_c21b49ee),
    .b(al_31a3e7af[211]),
    .c(al_955db046[211]),
    .o(al_b0408eb[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3e9bdfd0 (
    .a(al_c21b49ee),
    .b(al_31a3e7af[212]),
    .c(al_955db046[212]),
    .o(al_b0408eb[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c2bc58f (
    .a(al_c21b49ee),
    .b(al_31a3e7af[213]),
    .c(al_955db046[213]),
    .o(al_b0408eb[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_dffca741 (
    .a(al_c21b49ee),
    .b(al_31a3e7af[214]),
    .c(al_955db046[214]),
    .o(al_b0408eb[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7f2df993 (
    .a(al_c21b49ee),
    .b(al_31a3e7af[215]),
    .c(al_955db046[215]),
    .o(al_b0408eb[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9f58f555 (
    .a(al_b09bcab2),
    .b(al_31a3e7af[204]),
    .c(al_955db046[204]),
    .o(al_6b6ef69[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1491ea98 (
    .a(al_b09bcab2),
    .b(al_31a3e7af[205]),
    .c(al_955db046[205]),
    .o(al_6b6ef69[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b58a5cf1 (
    .a(al_b09bcab2),
    .b(al_31a3e7af[206]),
    .c(al_955db046[206]),
    .o(al_6b6ef69[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3cd69505 (
    .a(al_b09bcab2),
    .b(al_31a3e7af[207]),
    .c(al_955db046[207]),
    .o(al_6b6ef69[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a0990ad5 (
    .a(al_b09bcab2),
    .b(al_31a3e7af[208]),
    .c(al_955db046[208]),
    .o(al_6b6ef69[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_237ae028 (
    .a(al_b09bcab2),
    .b(al_31a3e7af[209]),
    .c(al_955db046[209]),
    .o(al_6b6ef69[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fa01ad0c (
    .a(al_b62a0a78),
    .b(al_31a3e7af[198]),
    .c(al_955db046[198]),
    .o(al_4c1bada4[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d46fdc0e (
    .a(al_b62a0a78),
    .b(al_31a3e7af[199]),
    .c(al_955db046[199]),
    .o(al_4c1bada4[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2ada342b (
    .a(al_b62a0a78),
    .b(al_31a3e7af[200]),
    .c(al_955db046[200]),
    .o(al_4c1bada4[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d6892319 (
    .a(al_b62a0a78),
    .b(al_31a3e7af[201]),
    .c(al_955db046[201]),
    .o(al_4c1bada4[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d5e1d07 (
    .a(al_b62a0a78),
    .b(al_31a3e7af[202]),
    .c(al_955db046[202]),
    .o(al_4c1bada4[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_506a8681 (
    .a(al_b62a0a78),
    .b(al_31a3e7af[203]),
    .c(al_955db046[203]),
    .o(al_4c1bada4[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b239d175 (
    .a(al_27d43db3),
    .b(al_31a3e7af[252]),
    .c(al_955db046[252]),
    .o(al_3ab36424[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a8573a5 (
    .a(al_27d43db3),
    .b(al_31a3e7af[253]),
    .c(al_955db046[253]),
    .o(al_3ab36424[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7772329e (
    .a(al_27d43db3),
    .b(al_31a3e7af[254]),
    .c(al_955db046[254]),
    .o(al_3ab36424[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_cf0aa803 (
    .a(al_27d43db3),
    .b(al_31a3e7af[255]),
    .c(al_955db046[255]),
    .o(al_3ab36424[3]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_e665a001 (
    .i(al_ee7571b0),
    .o(al_326d3b34[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9bc2d53c (
    .i(al_326d3b34[0]),
    .o(al_9a6187ef));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8a18c0a0 (
    .i(al_e6d4af1),
    .o(al_326d3b34[10]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_5bec2ce6 (
    .i(al_326d3b34[10]),
    .o(al_815c8034));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f185147f (
    .i(al_1759a3a0),
    .o(al_326d3b34[11]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_fcbc391c (
    .i(al_326d3b34[11]),
    .o(al_87f40037));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d4e775d6 (
    .i(al_30c9bd77),
    .o(al_326d3b34[12]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d709034b (
    .i(al_326d3b34[12]),
    .o(al_843f6bac));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4b7e59b9 (
    .i(al_6f07b96e),
    .o(al_326d3b34[13]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_dccb4aa7 (
    .i(al_326d3b34[13]),
    .o(al_535f72cd));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_91e78b5a (
    .i(al_4ab9f9ad),
    .o(al_326d3b34[14]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_edf92877 (
    .i(al_326d3b34[14]),
    .o(al_17b42586));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_170f9f54 (
    .i(al_7c6973e),
    .o(al_326d3b34[15]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b6cbfd02 (
    .i(al_326d3b34[15]),
    .o(al_df90085e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_fba949ff (
    .i(al_1f596d24),
    .o(al_326d3b34[16]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9a7310d3 (
    .i(al_326d3b34[16]),
    .o(al_72ab91cb));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d7f1343d (
    .i(al_dc57999f),
    .o(al_326d3b34[17]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4651e15 (
    .i(al_326d3b34[17]),
    .o(al_c9d182cf));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c9d1f4d6 (
    .i(al_f9e69b00),
    .o(al_326d3b34[18]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9c38be14 (
    .i(al_326d3b34[18]),
    .o(al_4f9aa153));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_45d5e5aa (
    .i(al_3a2d553d),
    .o(al_326d3b34[19]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_fd371e13 (
    .i(al_326d3b34[19]),
    .o(al_d4c409ba));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_aed312d6 (
    .i(al_b0c5cb0b),
    .o(al_326d3b34[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d8a34105 (
    .i(al_326d3b34[1]),
    .o(al_e2476620));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4cbdc0dd (
    .i(al_a88d3bd8),
    .o(al_326d3b34[20]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2a992704 (
    .i(al_326d3b34[20]),
    .o(al_24944e5c));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_75661408 (
    .i(al_722c0dcd),
    .o(al_326d3b34[21]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3f59adbd (
    .i(al_326d3b34[21]),
    .o(al_e2f3bed2));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_45f61156 (
    .i(al_4e018b61),
    .o(al_326d3b34[22]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_35ce69c6 (
    .i(al_326d3b34[22]),
    .o(al_6db10ea9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_63f89d75 (
    .i(al_1f414bbe),
    .o(al_326d3b34[23]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_17006966 (
    .i(al_326d3b34[23]),
    .o(al_7bbb36d3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3f473fdb (
    .i(al_eadb4e14),
    .o(al_326d3b34[24]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_17d0c151 (
    .i(al_326d3b34[24]),
    .o(al_8d8df5a3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f6433141 (
    .i(al_a771a309),
    .o(al_326d3b34[25]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c0034ebf (
    .i(al_326d3b34[25]),
    .o(al_2fc8b96e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5bcedd06 (
    .i(al_20f5f77c),
    .o(al_326d3b34[26]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_33e70645 (
    .i(al_326d3b34[26]),
    .o(al_d27a1279));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_bc09b63a (
    .i(al_d88aee38),
    .o(al_326d3b34[27]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d31abbe6 (
    .i(al_326d3b34[27]),
    .o(al_a48594d3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_eb8ff375 (
    .i(al_f9c30b23),
    .o(al_326d3b34[28]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_427cdee4 (
    .i(al_326d3b34[28]),
    .o(al_521fd670));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_14aa8090 (
    .i(al_d2a2bf32),
    .o(al_326d3b34[29]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_936564d5 (
    .i(al_326d3b34[29]),
    .o(al_1919cac5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8c48aa19 (
    .i(al_b09b809),
    .o(al_326d3b34[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_39945100 (
    .i(al_326d3b34[2]),
    .o(al_6e50ac65));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_cc8d66b9 (
    .i(al_c41fccfb),
    .o(al_326d3b34[30]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_fd445655 (
    .i(al_326d3b34[30]),
    .o(al_8dc56974));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c0d8657d (
    .i(al_91458dff),
    .o(al_326d3b34[31]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_5596dec0 (
    .i(al_326d3b34[31]),
    .o(al_8b05cae6));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3619c3e3 (
    .i(al_ade031de),
    .o(al_326d3b34[32]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c628c6d4 (
    .i(al_326d3b34[32]),
    .o(al_7bafa36d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_beb4aa7b (
    .i(al_830e948),
    .o(al_326d3b34[33]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c85f6968 (
    .i(al_326d3b34[33]),
    .o(al_25e4ab96));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_fd6dd438 (
    .i(al_d0276689),
    .o(al_326d3b34[34]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_54d77af1 (
    .i(al_326d3b34[34]),
    .o(al_6e370c03));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8fe3378a (
    .i(al_8e003744),
    .o(al_326d3b34[35]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d8becca1 (
    .i(al_326d3b34[35]),
    .o(al_770f9dd1));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ccc93ec9 (
    .i(al_8d08d03c),
    .o(al_326d3b34[36]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_163325e8 (
    .i(al_326d3b34[36]),
    .o(al_e2d4d651));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ddc39596 (
    .i(al_e470f61d),
    .o(al_326d3b34[37]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b9fc0d29 (
    .i(al_326d3b34[37]),
    .o(al_5be1fa83));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a50a5cfa (
    .i(al_93161d1e),
    .o(al_326d3b34[38]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_40f9f690 (
    .i(al_326d3b34[38]),
    .o(al_fd460907));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_cd3e9916 (
    .i(al_77d022d8),
    .o(al_326d3b34[39]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_248ac678 (
    .i(al_326d3b34[39]),
    .o(al_8815304a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ed69e41f (
    .i(al_ba71435f),
    .o(al_326d3b34[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_aeff1651 (
    .i(al_326d3b34[3]),
    .o(al_2e8aa91));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7181a51d (
    .i(al_c732c324),
    .o(al_326d3b34[40]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_17be58b7 (
    .i(al_326d3b34[40]),
    .o(al_ce1c71c5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_af4c071f (
    .i(al_fbdc3092),
    .o(al_326d3b34[41]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_33acf119 (
    .i(al_326d3b34[41]),
    .o(al_9929d21));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_625f87c2 (
    .i(al_142dd1c8),
    .o(al_326d3b34[42]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6faf0eb8 (
    .i(al_326d3b34[42]),
    .o(al_23ce284b));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c5995baf (
    .i(al_b40c9ab5),
    .o(al_326d3b34[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_642ddee6 (
    .i(al_326d3b34[4]),
    .o(al_4aba11ac));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1c4c81f0 (
    .i(al_fbbf0c04),
    .o(al_326d3b34[5]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e8f1fafb (
    .i(al_326d3b34[5]),
    .o(al_20c1f74d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_bac212df (
    .i(al_335c3c71),
    .o(al_326d3b34[6]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c1517d6a (
    .i(al_326d3b34[6]),
    .o(al_8fa72152));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b072e92f (
    .i(al_be14e3f3),
    .o(al_326d3b34[7]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7a0924f9 (
    .i(al_326d3b34[7]),
    .o(al_ea6ecc89));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_41f01f26 (
    .i(al_31cf7bc9),
    .o(al_326d3b34[8]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c243cf91 (
    .i(al_326d3b34[8]),
    .o(al_10f5be33));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3257cf24 (
    .i(al_8e660235),
    .o(al_326d3b34[9]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b009f188 (
    .i(al_326d3b34[9]),
    .o(al_d90f1fe1));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_df030cad (
    .a(al_37663fe4[0]),
    .b(al_37663fe4[1]),
    .c(al_37663fe4[2]),
    .d(al_37663fe4[3]),
    .e(al_37663fe4[4]),
    .f(al_7bafa36d),
    .o(al_852588b2));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_6f198553 (
    .a(al_d44a73a0[0]),
    .b(al_d44a73a0[1]),
    .c(al_d44a73a0[2]),
    .d(al_d44a73a0[3]),
    .e(al_d44a73a0[4]),
    .f(al_8b05cae6),
    .o(al_664e4e8f));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_864aae4d (
    .a(al_c244bf8b[0]),
    .b(al_c244bf8b[1]),
    .c(al_c244bf8b[2]),
    .d(al_c244bf8b[3]),
    .e(al_c244bf8b[4]),
    .f(al_8dc56974),
    .o(al_6f9c4eba));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_41401caf (
    .a(al_b04a4cbc[0]),
    .b(al_b04a4cbc[1]),
    .c(al_b04a4cbc[2]),
    .d(al_b04a4cbc[3]),
    .e(al_b04a4cbc[4]),
    .f(al_1919cac5),
    .o(al_55b9d73d));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_c407e023 (
    .a(al_ead25ba5[0]),
    .b(al_ead25ba5[1]),
    .c(al_ead25ba5[2]),
    .d(al_ead25ba5[3]),
    .e(al_ead25ba5[4]),
    .f(al_521fd670),
    .o(al_3858b210));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_26a79c5e (
    .a(al_206e4ef2[0]),
    .b(al_206e4ef2[1]),
    .c(al_206e4ef2[2]),
    .d(al_206e4ef2[3]),
    .e(al_206e4ef2[4]),
    .f(al_a48594d3),
    .o(al_96b7453));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_2ea505aa (
    .a(al_4f6bae56[0]),
    .b(al_4f6bae56[1]),
    .c(al_4f6bae56[2]),
    .d(al_4f6bae56[3]),
    .e(al_4f6bae56[4]),
    .f(al_d27a1279),
    .o(al_ee3904b1));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_68b86d88 (
    .a(al_5c6ba19f[0]),
    .b(al_5c6ba19f[1]),
    .c(al_5c6ba19f[2]),
    .d(al_5c6ba19f[3]),
    .e(al_5c6ba19f[4]),
    .f(al_2fc8b96e),
    .o(al_1abf75fc));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_13e06972 (
    .a(al_430dd919[0]),
    .b(al_430dd919[1]),
    .c(al_430dd919[2]),
    .d(al_430dd919[3]),
    .e(al_430dd919[4]),
    .f(al_8d8df5a3),
    .o(al_f9fd3044));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_f6ea2936 (
    .a(al_269b6545[0]),
    .b(al_269b6545[1]),
    .c(al_269b6545[2]),
    .d(al_269b6545[3]),
    .e(al_269b6545[4]),
    .f(al_7bbb36d3),
    .o(al_14656fdb));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_e25dfbac (
    .a(al_d9591ec3[0]),
    .b(al_d9591ec3[1]),
    .c(al_d9591ec3[2]),
    .d(al_d9591ec3[3]),
    .e(al_d9591ec3[4]),
    .f(al_9929d21),
    .o(al_7aee3607));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_2415086a (
    .a(al_384dd51d[0]),
    .b(al_384dd51d[1]),
    .c(al_384dd51d[2]),
    .d(al_384dd51d[3]),
    .e(al_384dd51d[4]),
    .f(al_6db10ea9),
    .o(al_130738c8));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_eb454ef9 (
    .a(al_55ef04c8[0]),
    .b(al_55ef04c8[1]),
    .c(al_55ef04c8[2]),
    .d(al_55ef04c8[3]),
    .e(al_55ef04c8[4]),
    .f(al_e2f3bed2),
    .o(al_f45ad02a));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_627f153f (
    .a(al_9cdd3a01[0]),
    .b(al_9cdd3a01[1]),
    .c(al_9cdd3a01[2]),
    .d(al_9cdd3a01[3]),
    .e(al_9cdd3a01[4]),
    .f(al_24944e5c),
    .o(al_4783da3f));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_a8f8db88 (
    .a(al_f5e6b3f5[0]),
    .b(al_f5e6b3f5[1]),
    .c(al_f5e6b3f5[2]),
    .d(al_f5e6b3f5[3]),
    .e(al_f5e6b3f5[4]),
    .f(al_d4c409ba),
    .o(al_b285e414));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_67e31978 (
    .a(al_175608a7[0]),
    .b(al_175608a7[1]),
    .c(al_175608a7[2]),
    .d(al_175608a7[3]),
    .e(al_175608a7[4]),
    .f(al_4f9aa153),
    .o(al_ef6d9f73));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_bb60c673 (
    .a(al_8af537d6[0]),
    .b(al_8af537d6[1]),
    .c(al_8af537d6[2]),
    .d(al_8af537d6[3]),
    .e(al_8af537d6[4]),
    .f(al_c9d182cf),
    .o(al_a7a585be));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_30b72b72 (
    .a(al_2d22d77a[0]),
    .b(al_2d22d77a[1]),
    .c(al_2d22d77a[2]),
    .d(al_2d22d77a[3]),
    .e(al_2d22d77a[4]),
    .f(al_72ab91cb),
    .o(al_3f68feff));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_1bd8fb12 (
    .a(al_100c2219[0]),
    .b(al_100c2219[1]),
    .c(al_100c2219[2]),
    .d(al_100c2219[3]),
    .e(al_100c2219[4]),
    .f(al_df90085e),
    .o(al_92250858));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_18942ff4 (
    .a(al_71242bdd[0]),
    .b(al_71242bdd[1]),
    .c(al_71242bdd[2]),
    .d(al_71242bdd[3]),
    .e(al_71242bdd[4]),
    .f(al_17b42586),
    .o(al_b4d25a49));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_d93aebaf (
    .a(al_44864e28[0]),
    .b(al_44864e28[1]),
    .c(al_44864e28[2]),
    .d(al_44864e28[3]),
    .e(al_44864e28[4]),
    .f(al_535f72cd),
    .o(al_3b280eeb));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_3355439 (
    .a(al_2119f32d[0]),
    .b(al_2119f32d[1]),
    .c(al_2119f32d[2]),
    .d(al_2119f32d[3]),
    .e(al_2119f32d[4]),
    .f(al_ce1c71c5),
    .o(al_cda79e31));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_f3786c72 (
    .a(al_4206b0c2[0]),
    .b(al_4206b0c2[1]),
    .c(al_4206b0c2[2]),
    .d(al_4206b0c2[3]),
    .e(al_4206b0c2[4]),
    .f(al_843f6bac),
    .o(al_a07095e8));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_b6287b90 (
    .a(al_d6b9e41[0]),
    .b(al_d6b9e41[1]),
    .c(al_d6b9e41[2]),
    .d(al_d6b9e41[3]),
    .e(al_d6b9e41[4]),
    .f(al_87f40037),
    .o(al_bf50c51c));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_61fd8b4b (
    .a(al_b5082a19[0]),
    .b(al_b5082a19[1]),
    .c(al_b5082a19[2]),
    .d(al_b5082a19[3]),
    .e(al_b5082a19[4]),
    .f(al_815c8034),
    .o(al_472a7b46));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_79145387 (
    .a(al_56e72bf4[0]),
    .b(al_56e72bf4[1]),
    .c(al_56e72bf4[2]),
    .d(al_56e72bf4[3]),
    .e(al_56e72bf4[4]),
    .f(al_d90f1fe1),
    .o(al_b9b495b9));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_9f7d9f4f (
    .a(al_46e8788c[0]),
    .b(al_46e8788c[1]),
    .c(al_46e8788c[2]),
    .d(al_46e8788c[3]),
    .e(al_46e8788c[4]),
    .f(al_10f5be33),
    .o(al_4531bc64));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_8160148 (
    .a(al_d61bccef[0]),
    .b(al_d61bccef[1]),
    .c(al_d61bccef[2]),
    .d(al_d61bccef[3]),
    .e(al_d61bccef[4]),
    .f(al_ea6ecc89),
    .o(al_3f7b50be));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_19a4f8d (
    .a(al_1e255230[0]),
    .b(al_1e255230[1]),
    .c(al_1e255230[2]),
    .d(al_1e255230[3]),
    .e(al_1e255230[4]),
    .f(al_8fa72152),
    .o(al_4cb605a3));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_2004527b (
    .a(al_d9be1f39[0]),
    .b(al_d9be1f39[1]),
    .c(al_d9be1f39[2]),
    .d(al_d9be1f39[3]),
    .e(al_d9be1f39[4]),
    .f(al_20c1f74d),
    .o(al_2ebef479));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_84f24aa5 (
    .a(al_f78383db[0]),
    .b(al_f78383db[1]),
    .c(al_f78383db[2]),
    .d(al_f78383db[3]),
    .e(al_f78383db[4]),
    .f(al_4aba11ac),
    .o(al_d93c50d7));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_6a4e1d29 (
    .a(al_4a30bd0f[0]),
    .b(al_4a30bd0f[1]),
    .c(al_4a30bd0f[2]),
    .d(al_4a30bd0f[3]),
    .e(al_4a30bd0f[4]),
    .f(al_2e8aa91),
    .o(al_6a0200a0));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_3aaef238 (
    .a(al_662b3089[0]),
    .b(al_662b3089[1]),
    .c(al_662b3089[2]),
    .d(al_662b3089[3]),
    .e(al_662b3089[4]),
    .f(al_8815304a),
    .o(al_e3bba389));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_c29e6a0b (
    .a(al_6b9e1d84[0]),
    .b(al_6b9e1d84[1]),
    .c(al_6b9e1d84[2]),
    .d(al_6b9e1d84[3]),
    .e(al_6b9e1d84[4]),
    .f(al_6e50ac65),
    .o(al_ce868614));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_14594dd2 (
    .a(al_abd25e4c[0]),
    .b(al_abd25e4c[1]),
    .c(al_abd25e4c[2]),
    .d(al_abd25e4c[3]),
    .e(al_abd25e4c[4]),
    .f(al_e2476620),
    .o(al_89b57934));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_6e4fedea (
    .a(al_5362aaf[0]),
    .b(al_5362aaf[1]),
    .c(al_5362aaf[2]),
    .d(al_5362aaf[3]),
    .e(al_5362aaf[4]),
    .f(al_9a6187ef),
    .o(al_d6502391));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_dd9ba371 (
    .a(al_2ef171e7[0]),
    .b(al_2ef171e7[1]),
    .c(al_2ef171e7[2]),
    .d(al_2ef171e7[3]),
    .e(al_2ef171e7[4]),
    .f(al_fd460907),
    .o(al_15554a76));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_4b81127f (
    .a(al_8349e0d1[0]),
    .b(al_8349e0d1[1]),
    .c(al_8349e0d1[2]),
    .d(al_8349e0d1[3]),
    .e(al_8349e0d1[4]),
    .f(al_5be1fa83),
    .o(al_b57594f0));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_73da5792 (
    .a(al_e31889d8[0]),
    .b(al_e31889d8[1]),
    .c(al_e31889d8[2]),
    .d(al_e31889d8[3]),
    .e(al_e31889d8[4]),
    .f(al_e2d4d651),
    .o(al_ca5b293f));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_185ad957 (
    .a(al_85a14e36[0]),
    .b(al_85a14e36[1]),
    .c(al_85a14e36[2]),
    .d(al_85a14e36[3]),
    .e(al_85a14e36[4]),
    .f(al_770f9dd1),
    .o(al_da329b96));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_4a3a1b20 (
    .a(al_f359f0c8[0]),
    .b(al_f359f0c8[1]),
    .c(al_f359f0c8[2]),
    .d(al_f359f0c8[3]),
    .e(al_f359f0c8[4]),
    .f(al_6e370c03),
    .o(al_f3b50940));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_4b1a6527 (
    .a(al_e865b87a[0]),
    .b(al_e865b87a[1]),
    .c(al_e865b87a[2]),
    .d(al_e865b87a[3]),
    .e(al_e865b87a[4]),
    .f(al_25e4ab96),
    .o(al_14200974));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_f6e3fbac (
    .a(al_1d102248[0]),
    .b(al_1d102248[1]),
    .c(al_1d102248[2]),
    .d(al_1d102248[3]),
    .e(al_1d102248[4]),
    .f(al_23ce284b),
    .o(al_d9a683f3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b2dd6461 (
    .i(al_4cc6df6e),
    .o(al_57f9dbc3[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_eb7117ba (
    .i(al_57f9dbc3[0]),
    .o(al_b8212fd4));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_5d55d84a (
    .a(al_99c75e01),
    .b(al_9a6187ef),
    .o(al_4cc6df6e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d39cf9d1 (
    .i(al_cae86888),
    .o(al_57f9dbc3[10]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_40f50d78 (
    .i(al_57f9dbc3[10]),
    .o(al_1584b2ff));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_d9e513c2 (
    .a(al_99c75e01),
    .b(al_815c8034),
    .o(al_cae86888));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4fed4911 (
    .i(al_db0962eb),
    .o(al_57f9dbc3[11]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a2814582 (
    .i(al_57f9dbc3[11]),
    .o(al_e463a453));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_658c66f3 (
    .a(al_99c75e01),
    .b(al_87f40037),
    .o(al_db0962eb));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5b30d4da (
    .i(al_4d350d21),
    .o(al_57f9dbc3[12]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_26d975a0 (
    .i(al_57f9dbc3[12]),
    .o(al_952b0ccf));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_28b765f4 (
    .a(al_99c75e01),
    .b(al_843f6bac),
    .o(al_4d350d21));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7f584982 (
    .i(al_925b7c77),
    .o(al_57f9dbc3[13]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1922130f (
    .i(al_57f9dbc3[13]),
    .o(al_bf72b0fb));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_fe9ea46d (
    .a(al_99c75e01),
    .b(al_535f72cd),
    .o(al_925b7c77));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_cf1b46a2 (
    .i(al_f8edc4ff),
    .o(al_57f9dbc3[14]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_cd0475 (
    .i(al_57f9dbc3[14]),
    .o(al_221290fc));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_54ab92e1 (
    .a(al_99c75e01),
    .b(al_17b42586),
    .o(al_f8edc4ff));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_478bd8a9 (
    .i(al_77720e8a),
    .o(al_57f9dbc3[15]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1a67ff78 (
    .i(al_57f9dbc3[15]),
    .o(al_fd118264));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_6430637e (
    .a(al_99c75e01),
    .b(al_df90085e),
    .o(al_77720e8a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_be704e59 (
    .i(al_556566a0),
    .o(al_57f9dbc3[16]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_f0df58de (
    .i(al_57f9dbc3[16]),
    .o(al_f3b3330));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_2eefdac4 (
    .a(al_99c75e01),
    .b(al_72ab91cb),
    .o(al_556566a0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4f142844 (
    .i(al_69a4bab5),
    .o(al_57f9dbc3[17]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4b0051c4 (
    .i(al_57f9dbc3[17]),
    .o(al_6adcd3f0));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_50c8bedd (
    .a(al_99c75e01),
    .b(al_c9d182cf),
    .o(al_69a4bab5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_cc720022 (
    .i(al_db74407e),
    .o(al_57f9dbc3[18]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_19ffb72 (
    .i(al_57f9dbc3[18]),
    .o(al_dd36eaa4));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_dd6e9b7b (
    .a(al_99c75e01),
    .b(al_4f9aa153),
    .o(al_db74407e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3c4cfcce (
    .i(al_787c471e),
    .o(al_57f9dbc3[19]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c48f5d82 (
    .i(al_57f9dbc3[19]),
    .o(al_7c446883));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_12f848c7 (
    .a(al_99c75e01),
    .b(al_d4c409ba),
    .o(al_787c471e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3f747b75 (
    .i(al_1e064d5f),
    .o(al_57f9dbc3[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_421b5b13 (
    .i(al_57f9dbc3[1]),
    .o(al_86df7d12));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_edbb1ac2 (
    .a(al_99c75e01),
    .b(al_e2476620),
    .o(al_1e064d5f));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ca2958f6 (
    .i(al_c03f902b),
    .o(al_57f9dbc3[20]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9b056c87 (
    .i(al_57f9dbc3[20]),
    .o(al_1591047a));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_1d4b8950 (
    .a(al_99c75e01),
    .b(al_24944e5c),
    .o(al_c03f902b));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_794ddfd9 (
    .i(al_3e851499),
    .o(al_57f9dbc3[21]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_f208b289 (
    .i(al_57f9dbc3[21]),
    .o(al_d3c4d360));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_5366f82f (
    .a(al_99c75e01),
    .b(al_e2f3bed2),
    .o(al_3e851499));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1daffa2a (
    .i(al_6652ce21),
    .o(al_57f9dbc3[22]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6e8a79a8 (
    .i(al_57f9dbc3[22]),
    .o(al_6d6760dd));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_85bc2e2 (
    .a(al_99c75e01),
    .b(al_6db10ea9),
    .o(al_6652ce21));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7709cb3f (
    .i(al_4f8f3ec),
    .o(al_57f9dbc3[23]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_46defc19 (
    .i(al_57f9dbc3[23]),
    .o(al_9cf6a965));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_27ce07d1 (
    .a(al_99c75e01),
    .b(al_7bbb36d3),
    .o(al_4f8f3ec));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_557daaa5 (
    .i(al_5b5189ed),
    .o(al_57f9dbc3[24]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c32e1b48 (
    .i(al_57f9dbc3[24]),
    .o(al_37a8c4a3));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_b24d776 (
    .a(al_99c75e01),
    .b(al_8d8df5a3),
    .o(al_5b5189ed));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b72701a0 (
    .i(al_92cbdd49),
    .o(al_57f9dbc3[25]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_664301d3 (
    .i(al_57f9dbc3[25]),
    .o(al_2c31bcd7));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_e6ffb830 (
    .a(al_99c75e01),
    .b(al_2fc8b96e),
    .o(al_92cbdd49));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c1950e (
    .i(al_d55891ef),
    .o(al_57f9dbc3[26]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_230f7ffb (
    .i(al_57f9dbc3[26]),
    .o(al_bbe31482));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_8db7dbc0 (
    .a(al_99c75e01),
    .b(al_d27a1279),
    .o(al_d55891ef));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7a0e27f6 (
    .i(al_ef98f3e9),
    .o(al_57f9dbc3[27]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_eb997022 (
    .i(al_57f9dbc3[27]),
    .o(al_edff11e6));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_651b7a8 (
    .a(al_99c75e01),
    .b(al_a48594d3),
    .o(al_ef98f3e9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c01e8220 (
    .i(al_1c0f25b0),
    .o(al_57f9dbc3[28]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_af88d0f5 (
    .i(al_57f9dbc3[28]),
    .o(al_4b287773));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_12d2f49b (
    .a(al_99c75e01),
    .b(al_521fd670),
    .o(al_1c0f25b0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_40083931 (
    .i(al_70ff6ecf),
    .o(al_57f9dbc3[29]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_dfb045db (
    .i(al_57f9dbc3[29]),
    .o(al_a18a78ec));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_d40e521f (
    .a(al_99c75e01),
    .b(al_1919cac5),
    .o(al_70ff6ecf));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_6523a7fe (
    .i(al_deb7c4e9),
    .o(al_57f9dbc3[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7d267a91 (
    .i(al_57f9dbc3[2]),
    .o(al_f8b11b95));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_9b7064ac (
    .a(al_99c75e01),
    .b(al_6e50ac65),
    .o(al_deb7c4e9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_df29deb9 (
    .i(al_a0a92d29),
    .o(al_57f9dbc3[30]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_602ec6ed (
    .i(al_57f9dbc3[30]),
    .o(al_dd0c66b3));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_adf63227 (
    .a(al_99c75e01),
    .b(al_8dc56974),
    .o(al_a0a92d29));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_cd7dc5c3 (
    .i(al_dc8a13dc),
    .o(al_57f9dbc3[31]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_deed8d4b (
    .i(al_57f9dbc3[31]),
    .o(al_edb83574));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_26650a51 (
    .a(al_99c75e01),
    .b(al_8b05cae6),
    .o(al_dc8a13dc));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_51f1f78 (
    .i(al_41f57e5d),
    .o(al_57f9dbc3[32]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_706a57ab (
    .i(al_57f9dbc3[32]),
    .o(al_2935d0ed));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_3c388017 (
    .a(al_99c75e01),
    .b(al_7bafa36d),
    .o(al_41f57e5d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_e8f765df (
    .i(al_b3610ba2),
    .o(al_57f9dbc3[33]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_65ec8102 (
    .i(al_57f9dbc3[33]),
    .o(al_538eda90));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_f7da6e9 (
    .a(al_99c75e01),
    .b(al_25e4ab96),
    .o(al_b3610ba2));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_532f7ae6 (
    .i(al_95dd6731),
    .o(al_57f9dbc3[34]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7e01eec3 (
    .i(al_57f9dbc3[34]),
    .o(al_2503fdb));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_6b4abe8d (
    .a(al_99c75e01),
    .b(al_6e370c03),
    .o(al_95dd6731));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_39dff613 (
    .i(al_9f893f0c),
    .o(al_57f9dbc3[35]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_cf5284f2 (
    .i(al_57f9dbc3[35]),
    .o(al_f8fcd204));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_fbc705c1 (
    .a(al_99c75e01),
    .b(al_770f9dd1),
    .o(al_9f893f0c));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_2a9eee20 (
    .i(al_8ad430a7),
    .o(al_57f9dbc3[36]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2aedde8e (
    .i(al_57f9dbc3[36]),
    .o(al_467a2ca));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_1cfba62 (
    .a(al_99c75e01),
    .b(al_e2d4d651),
    .o(al_8ad430a7));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_2b43fc58 (
    .i(al_c446e1c1),
    .o(al_57f9dbc3[37]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_cbf2a181 (
    .i(al_57f9dbc3[37]),
    .o(al_c76ae5c3));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_f4282fec (
    .a(al_99c75e01),
    .b(al_5be1fa83),
    .o(al_c446e1c1));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4b81515a (
    .i(al_ec12476e),
    .o(al_57f9dbc3[38]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6ac9aa43 (
    .i(al_57f9dbc3[38]),
    .o(al_d2c8f1b1));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_c599b309 (
    .a(al_99c75e01),
    .b(al_fd460907),
    .o(al_ec12476e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_86262675 (
    .i(al_1a61307),
    .o(al_57f9dbc3[39]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_5ae895a3 (
    .i(al_57f9dbc3[39]),
    .o(al_282d371d));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_b2fedee4 (
    .a(al_99c75e01),
    .b(al_8815304a),
    .o(al_1a61307));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_fa42d09c (
    .i(al_199f1a83),
    .o(al_57f9dbc3[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_44e0b84c (
    .i(al_57f9dbc3[3]),
    .o(al_cd27f05c));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_e7ce22b6 (
    .a(al_99c75e01),
    .b(al_2e8aa91),
    .o(al_199f1a83));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b9824160 (
    .i(al_a04a63e0),
    .o(al_57f9dbc3[40]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_cf3e5351 (
    .i(al_57f9dbc3[40]),
    .o(al_27b77d58));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_9406b689 (
    .a(al_99c75e01),
    .b(al_ce1c71c5),
    .o(al_a04a63e0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_18fb7f52 (
    .i(al_2a05599e),
    .o(al_57f9dbc3[41]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_dcff7ae1 (
    .i(al_57f9dbc3[41]),
    .o(al_d4d145cc));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_191e03f8 (
    .a(al_99c75e01),
    .b(al_9929d21),
    .o(al_2a05599e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_67bf5cfa (
    .i(al_61d4d1dd),
    .o(al_57f9dbc3[42]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_83675ce1 (
    .i(al_57f9dbc3[42]),
    .o(al_129a2529));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_5231d2c7 (
    .a(al_99c75e01),
    .b(al_23ce284b),
    .o(al_61d4d1dd));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_187c0b35 (
    .i(al_bcb98901),
    .o(al_57f9dbc3[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_36baad26 (
    .i(al_57f9dbc3[4]),
    .o(al_14cefac2));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_8ff2053a (
    .a(al_99c75e01),
    .b(al_4aba11ac),
    .o(al_bcb98901));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4f3cbea1 (
    .i(al_3c6c8ee5),
    .o(al_57f9dbc3[5]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b7bbef60 (
    .i(al_57f9dbc3[5]),
    .o(al_6fd6ffff));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_324f4c9e (
    .a(al_99c75e01),
    .b(al_20c1f74d),
    .o(al_3c6c8ee5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_26d0ab (
    .i(al_a1041e9),
    .o(al_57f9dbc3[6]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7ce690c1 (
    .i(al_57f9dbc3[6]),
    .o(al_f645b571));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_73877c82 (
    .a(al_99c75e01),
    .b(al_8fa72152),
    .o(al_a1041e9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b7f6b909 (
    .i(al_6bd0f993),
    .o(al_57f9dbc3[7]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d9496f7e (
    .i(al_57f9dbc3[7]),
    .o(al_3419432c));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_415d525a (
    .a(al_99c75e01),
    .b(al_ea6ecc89),
    .o(al_6bd0f993));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8218abb (
    .i(al_e0c544fc),
    .o(al_57f9dbc3[8]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7c4d708d (
    .i(al_57f9dbc3[8]),
    .o(al_b9e4ee74));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_74ebcf44 (
    .a(al_99c75e01),
    .b(al_10f5be33),
    .o(al_e0c544fc));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f077445e (
    .i(al_e5334d53),
    .o(al_57f9dbc3[9]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_951c70ab (
    .i(al_57f9dbc3[9]),
    .o(al_4b747cba));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_20f95737 (
    .a(al_99c75e01),
    .b(al_d90f1fe1),
    .o(al_e5334d53));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_8666cdcf (
    .a(al_5362aaf[0]),
    .b(al_4b4a698a),
    .o(al_aa09a9e5[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_84cc7655 (
    .a(al_5362aaf[0]),
    .b(al_5362aaf[1]),
    .c(al_4b4a698a),
    .o(al_aa09a9e5[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_ec20055e (
    .a(al_5362aaf[0]),
    .b(al_5362aaf[1]),
    .c(al_5362aaf[2]),
    .d(al_4b4a698a),
    .o(al_aa09a9e5[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_64c90d4a (
    .a(al_5362aaf[0]),
    .b(al_5362aaf[1]),
    .c(al_5362aaf[2]),
    .d(al_5362aaf[3]),
    .e(al_4b4a698a),
    .o(al_aa09a9e5[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_9d4e3f92 (
    .a(al_5362aaf[0]),
    .b(al_5362aaf[1]),
    .c(al_5362aaf[2]),
    .d(al_5362aaf[3]),
    .e(al_5362aaf[4]),
    .f(al_4b4a698a),
    .o(al_aa09a9e5[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2d3ace4 (
    .di(al_31a3e7af[5:4]),
    .raddr(al_aa09a9e5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_b8212fd4),
    .rdo(al_955db046[5:4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2b83018 (
    .di(al_31a3e7af[3:2]),
    .raddr(al_aa09a9e5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_b8212fd4),
    .rdo(al_955db046[3:2]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_73a0a39 (
    .di(al_31a3e7af[1:0]),
    .raddr(al_aa09a9e5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_b8212fd4),
    .rdo(al_955db046[1:0]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_4c119cf5 (
    .a(al_b5082a19[0]),
    .b(al_b8cc00cf),
    .o(al_4c8ce587[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_5fe2bf96 (
    .a(al_b5082a19[0]),
    .b(al_b5082a19[1]),
    .c(al_b8cc00cf),
    .o(al_4c8ce587[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_e9eb5c61 (
    .a(al_b5082a19[0]),
    .b(al_b5082a19[1]),
    .c(al_b5082a19[2]),
    .d(al_b8cc00cf),
    .o(al_4c8ce587[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_29756156 (
    .a(al_b5082a19[0]),
    .b(al_b5082a19[1]),
    .c(al_b5082a19[2]),
    .d(al_b5082a19[3]),
    .e(al_b8cc00cf),
    .o(al_4c8ce587[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_d545ac9a (
    .a(al_b5082a19[0]),
    .b(al_b5082a19[1]),
    .c(al_b5082a19[2]),
    .d(al_b5082a19[3]),
    .e(al_b5082a19[4]),
    .f(al_b8cc00cf),
    .o(al_4c8ce587[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9d2220ef (
    .di(al_31a3e7af[65:64]),
    .raddr(al_4c8ce587),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_1584b2ff),
    .rdo(al_955db046[65:64]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b8a1757 (
    .di(al_31a3e7af[63:62]),
    .raddr(al_4c8ce587),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_1584b2ff),
    .rdo(al_955db046[63:62]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b6d00bf5 (
    .di(al_31a3e7af[61:60]),
    .raddr(al_4c8ce587),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_1584b2ff),
    .rdo(al_955db046[61:60]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_a156315b (
    .a(al_d6b9e41[0]),
    .b(al_106fddab),
    .o(al_3854534a[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_3b9d61f1 (
    .a(al_d6b9e41[0]),
    .b(al_d6b9e41[1]),
    .c(al_106fddab),
    .o(al_3854534a[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_7cea5f1b (
    .a(al_d6b9e41[0]),
    .b(al_d6b9e41[1]),
    .c(al_d6b9e41[2]),
    .d(al_106fddab),
    .o(al_3854534a[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_5176d61 (
    .a(al_d6b9e41[0]),
    .b(al_d6b9e41[1]),
    .c(al_d6b9e41[2]),
    .d(al_d6b9e41[3]),
    .e(al_106fddab),
    .o(al_3854534a[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_a9937a5e (
    .a(al_d6b9e41[0]),
    .b(al_d6b9e41[1]),
    .c(al_d6b9e41[2]),
    .d(al_d6b9e41[3]),
    .e(al_d6b9e41[4]),
    .f(al_106fddab),
    .o(al_3854534a[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ef4dd470 (
    .di(al_31a3e7af[71:70]),
    .raddr(al_3854534a),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_e463a453),
    .rdo(al_955db046[71:70]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_fb5ad7cc (
    .di(al_31a3e7af[69:68]),
    .raddr(al_3854534a),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_e463a453),
    .rdo(al_955db046[69:68]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c52d3ed4 (
    .di(al_31a3e7af[67:66]),
    .raddr(al_3854534a),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_e463a453),
    .rdo(al_955db046[67:66]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_a7e98178 (
    .a(al_4206b0c2[0]),
    .b(al_82133c54),
    .o(al_49eb8970[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_c8df2a48 (
    .a(al_4206b0c2[0]),
    .b(al_4206b0c2[1]),
    .c(al_82133c54),
    .o(al_49eb8970[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_15c7cfd2 (
    .a(al_4206b0c2[0]),
    .b(al_4206b0c2[1]),
    .c(al_4206b0c2[2]),
    .d(al_82133c54),
    .o(al_49eb8970[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_f159dc0f (
    .a(al_4206b0c2[0]),
    .b(al_4206b0c2[1]),
    .c(al_4206b0c2[2]),
    .d(al_4206b0c2[3]),
    .e(al_82133c54),
    .o(al_49eb8970[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_4fa0887e (
    .a(al_4206b0c2[0]),
    .b(al_4206b0c2[1]),
    .c(al_4206b0c2[2]),
    .d(al_4206b0c2[3]),
    .e(al_4206b0c2[4]),
    .f(al_82133c54),
    .o(al_49eb8970[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_a56f4935 (
    .di(al_31a3e7af[77:76]),
    .raddr(al_49eb8970),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_952b0ccf),
    .rdo(al_955db046[77:76]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bdd55f5b (
    .di(al_31a3e7af[75:74]),
    .raddr(al_49eb8970),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_952b0ccf),
    .rdo(al_955db046[75:74]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_cd194947 (
    .di(al_31a3e7af[73:72]),
    .raddr(al_49eb8970),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_952b0ccf),
    .rdo(al_955db046[73:72]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_b4494c73 (
    .a(al_44864e28[0]),
    .b(al_9f6750b6),
    .o(al_39c7f0b5[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_832f32c2 (
    .a(al_44864e28[0]),
    .b(al_44864e28[1]),
    .c(al_9f6750b6),
    .o(al_39c7f0b5[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_50f9d5cd (
    .a(al_44864e28[0]),
    .b(al_44864e28[1]),
    .c(al_44864e28[2]),
    .d(al_9f6750b6),
    .o(al_39c7f0b5[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_52b309e3 (
    .a(al_44864e28[0]),
    .b(al_44864e28[1]),
    .c(al_44864e28[2]),
    .d(al_44864e28[3]),
    .e(al_9f6750b6),
    .o(al_39c7f0b5[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_a9e3c456 (
    .a(al_44864e28[0]),
    .b(al_44864e28[1]),
    .c(al_44864e28[2]),
    .d(al_44864e28[3]),
    .e(al_44864e28[4]),
    .f(al_9f6750b6),
    .o(al_39c7f0b5[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_645da486 (
    .di(al_31a3e7af[83:82]),
    .raddr(al_39c7f0b5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_bf72b0fb),
    .rdo(al_955db046[83:82]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_db66de46 (
    .di(al_31a3e7af[81:80]),
    .raddr(al_39c7f0b5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_bf72b0fb),
    .rdo(al_955db046[81:80]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_538b6f5 (
    .di(al_31a3e7af[79:78]),
    .raddr(al_39c7f0b5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_bf72b0fb),
    .rdo(al_955db046[79:78]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_1ae806ae (
    .a(al_71242bdd[0]),
    .b(al_21d51e65),
    .o(al_886fd669[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_7360c265 (
    .a(al_71242bdd[0]),
    .b(al_71242bdd[1]),
    .c(al_21d51e65),
    .o(al_886fd669[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_ccf03ebb (
    .a(al_71242bdd[0]),
    .b(al_71242bdd[1]),
    .c(al_71242bdd[2]),
    .d(al_21d51e65),
    .o(al_886fd669[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_bb5eea7 (
    .a(al_71242bdd[0]),
    .b(al_71242bdd[1]),
    .c(al_71242bdd[2]),
    .d(al_71242bdd[3]),
    .e(al_21d51e65),
    .o(al_886fd669[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_fba14472 (
    .a(al_71242bdd[0]),
    .b(al_71242bdd[1]),
    .c(al_71242bdd[2]),
    .d(al_71242bdd[3]),
    .e(al_71242bdd[4]),
    .f(al_21d51e65),
    .o(al_886fd669[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_5bb7b24f (
    .di(al_31a3e7af[89:88]),
    .raddr(al_886fd669),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_221290fc),
    .rdo(al_955db046[89:88]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3303b85c (
    .di(al_31a3e7af[87:86]),
    .raddr(al_886fd669),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_221290fc),
    .rdo(al_955db046[87:86]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_59287421 (
    .di(al_31a3e7af[85:84]),
    .raddr(al_886fd669),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_221290fc),
    .rdo(al_955db046[85:84]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_3668600b (
    .a(al_100c2219[0]),
    .b(al_3da9562a),
    .o(al_3550db07[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_32202c10 (
    .a(al_100c2219[0]),
    .b(al_100c2219[1]),
    .c(al_3da9562a),
    .o(al_3550db07[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_35cba2ca (
    .a(al_100c2219[0]),
    .b(al_100c2219[1]),
    .c(al_100c2219[2]),
    .d(al_3da9562a),
    .o(al_3550db07[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_33d064e2 (
    .a(al_100c2219[0]),
    .b(al_100c2219[1]),
    .c(al_100c2219[2]),
    .d(al_100c2219[3]),
    .e(al_3da9562a),
    .o(al_3550db07[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_5e7da843 (
    .a(al_100c2219[0]),
    .b(al_100c2219[1]),
    .c(al_100c2219[2]),
    .d(al_100c2219[3]),
    .e(al_100c2219[4]),
    .f(al_3da9562a),
    .o(al_3550db07[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_78f24769 (
    .di(al_31a3e7af[95:94]),
    .raddr(al_3550db07),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_fd118264),
    .rdo(al_955db046[95:94]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_cd9ff67c (
    .di(al_31a3e7af[93:92]),
    .raddr(al_3550db07),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_fd118264),
    .rdo(al_955db046[93:92]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_12818a28 (
    .di(al_31a3e7af[91:90]),
    .raddr(al_3550db07),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_fd118264),
    .rdo(al_955db046[91:90]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_3cd5b9f0 (
    .a(al_2d22d77a[0]),
    .b(al_d9d76d0a),
    .o(al_9823c42b[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_ff5ce183 (
    .a(al_2d22d77a[0]),
    .b(al_2d22d77a[1]),
    .c(al_d9d76d0a),
    .o(al_9823c42b[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_534ea3cb (
    .a(al_2d22d77a[0]),
    .b(al_2d22d77a[1]),
    .c(al_2d22d77a[2]),
    .d(al_d9d76d0a),
    .o(al_9823c42b[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_99541a12 (
    .a(al_2d22d77a[0]),
    .b(al_2d22d77a[1]),
    .c(al_2d22d77a[2]),
    .d(al_2d22d77a[3]),
    .e(al_d9d76d0a),
    .o(al_9823c42b[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_4c242a9 (
    .a(al_2d22d77a[0]),
    .b(al_2d22d77a[1]),
    .c(al_2d22d77a[2]),
    .d(al_2d22d77a[3]),
    .e(al_2d22d77a[4]),
    .f(al_d9d76d0a),
    .o(al_9823c42b[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_af927176 (
    .di(al_31a3e7af[101:100]),
    .raddr(al_9823c42b),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f3b3330),
    .rdo(al_955db046[101:100]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d288bb00 (
    .di(al_31a3e7af[99:98]),
    .raddr(al_9823c42b),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f3b3330),
    .rdo(al_955db046[99:98]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2d12520b (
    .di(al_31a3e7af[97:96]),
    .raddr(al_9823c42b),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f3b3330),
    .rdo(al_955db046[97:96]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e7afef21 (
    .a(al_8af537d6[0]),
    .b(al_64f79045),
    .o(al_90b3a908[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_cf87d06a (
    .a(al_8af537d6[0]),
    .b(al_8af537d6[1]),
    .c(al_64f79045),
    .o(al_90b3a908[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_bb934809 (
    .a(al_8af537d6[0]),
    .b(al_8af537d6[1]),
    .c(al_8af537d6[2]),
    .d(al_64f79045),
    .o(al_90b3a908[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_7a425a10 (
    .a(al_8af537d6[0]),
    .b(al_8af537d6[1]),
    .c(al_8af537d6[2]),
    .d(al_8af537d6[3]),
    .e(al_64f79045),
    .o(al_90b3a908[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_c983e1ac (
    .a(al_8af537d6[0]),
    .b(al_8af537d6[1]),
    .c(al_8af537d6[2]),
    .d(al_8af537d6[3]),
    .e(al_8af537d6[4]),
    .f(al_64f79045),
    .o(al_90b3a908[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_765a2290 (
    .di(al_31a3e7af[107:106]),
    .raddr(al_90b3a908),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6adcd3f0),
    .rdo(al_955db046[107:106]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e7a3e804 (
    .di(al_31a3e7af[105:104]),
    .raddr(al_90b3a908),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6adcd3f0),
    .rdo(al_955db046[105:104]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b5edc190 (
    .di(al_31a3e7af[103:102]),
    .raddr(al_90b3a908),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6adcd3f0),
    .rdo(al_955db046[103:102]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_45aa1448 (
    .a(al_175608a7[0]),
    .b(al_ab1b2b16),
    .o(al_61edc911[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_2495c760 (
    .a(al_175608a7[0]),
    .b(al_175608a7[1]),
    .c(al_ab1b2b16),
    .o(al_61edc911[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_2af8458a (
    .a(al_175608a7[0]),
    .b(al_175608a7[1]),
    .c(al_175608a7[2]),
    .d(al_ab1b2b16),
    .o(al_61edc911[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_daa2b9a6 (
    .a(al_175608a7[0]),
    .b(al_175608a7[1]),
    .c(al_175608a7[2]),
    .d(al_175608a7[3]),
    .e(al_ab1b2b16),
    .o(al_61edc911[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_c5e27616 (
    .a(al_175608a7[0]),
    .b(al_175608a7[1]),
    .c(al_175608a7[2]),
    .d(al_175608a7[3]),
    .e(al_175608a7[4]),
    .f(al_ab1b2b16),
    .o(al_61edc911[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7c663a0c (
    .di(al_31a3e7af[113:112]),
    .raddr(al_61edc911),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_dd36eaa4),
    .rdo(al_955db046[113:112]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_93495d83 (
    .di(al_31a3e7af[111:110]),
    .raddr(al_61edc911),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_dd36eaa4),
    .rdo(al_955db046[111:110]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_8f85f4c8 (
    .di(al_31a3e7af[109:108]),
    .raddr(al_61edc911),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_dd36eaa4),
    .rdo(al_955db046[109:108]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_9929a3a8 (
    .a(al_f5e6b3f5[0]),
    .b(al_c81182c),
    .o(al_abb88584[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_c5dd1c05 (
    .a(al_f5e6b3f5[0]),
    .b(al_f5e6b3f5[1]),
    .c(al_c81182c),
    .o(al_abb88584[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_88dd2f94 (
    .a(al_f5e6b3f5[0]),
    .b(al_f5e6b3f5[1]),
    .c(al_f5e6b3f5[2]),
    .d(al_c81182c),
    .o(al_abb88584[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_28b0b0fb (
    .a(al_f5e6b3f5[0]),
    .b(al_f5e6b3f5[1]),
    .c(al_f5e6b3f5[2]),
    .d(al_f5e6b3f5[3]),
    .e(al_c81182c),
    .o(al_abb88584[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_8b0efe0a (
    .a(al_f5e6b3f5[0]),
    .b(al_f5e6b3f5[1]),
    .c(al_f5e6b3f5[2]),
    .d(al_f5e6b3f5[3]),
    .e(al_f5e6b3f5[4]),
    .f(al_c81182c),
    .o(al_abb88584[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b16bac8d (
    .di(al_31a3e7af[119:118]),
    .raddr(al_abb88584),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_7c446883),
    .rdo(al_955db046[119:118]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_adb359fd (
    .di(al_31a3e7af[117:116]),
    .raddr(al_abb88584),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_7c446883),
    .rdo(al_955db046[117:116]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_82e1801 (
    .di(al_31a3e7af[115:114]),
    .raddr(al_abb88584),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_7c446883),
    .rdo(al_955db046[115:114]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_2c10e54 (
    .a(al_abd25e4c[0]),
    .b(al_9b5a4dbd),
    .o(al_3fe9a5bb[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_9c86265e (
    .a(al_abd25e4c[0]),
    .b(al_abd25e4c[1]),
    .c(al_9b5a4dbd),
    .o(al_3fe9a5bb[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_871a951a (
    .a(al_abd25e4c[0]),
    .b(al_abd25e4c[1]),
    .c(al_abd25e4c[2]),
    .d(al_9b5a4dbd),
    .o(al_3fe9a5bb[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_39053a64 (
    .a(al_abd25e4c[0]),
    .b(al_abd25e4c[1]),
    .c(al_abd25e4c[2]),
    .d(al_abd25e4c[3]),
    .e(al_9b5a4dbd),
    .o(al_3fe9a5bb[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_b97ecfb2 (
    .a(al_abd25e4c[0]),
    .b(al_abd25e4c[1]),
    .c(al_abd25e4c[2]),
    .d(al_abd25e4c[3]),
    .e(al_abd25e4c[4]),
    .f(al_9b5a4dbd),
    .o(al_3fe9a5bb[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f05156be (
    .di(al_31a3e7af[11:10]),
    .raddr(al_3fe9a5bb),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_86df7d12),
    .rdo(al_955db046[11:10]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bed2b77f (
    .di(al_31a3e7af[9:8]),
    .raddr(al_3fe9a5bb),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_86df7d12),
    .rdo(al_955db046[9:8]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_66646672 (
    .di(al_31a3e7af[7:6]),
    .raddr(al_3fe9a5bb),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_86df7d12),
    .rdo(al_955db046[7:6]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_5814326b (
    .a(al_9cdd3a01[0]),
    .b(al_b8da0e9e),
    .o(al_e94a3a72[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_dc4f9dbc (
    .a(al_9cdd3a01[0]),
    .b(al_9cdd3a01[1]),
    .c(al_b8da0e9e),
    .o(al_e94a3a72[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_a26d97f3 (
    .a(al_9cdd3a01[0]),
    .b(al_9cdd3a01[1]),
    .c(al_9cdd3a01[2]),
    .d(al_b8da0e9e),
    .o(al_e94a3a72[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_3ac6a3e1 (
    .a(al_9cdd3a01[0]),
    .b(al_9cdd3a01[1]),
    .c(al_9cdd3a01[2]),
    .d(al_9cdd3a01[3]),
    .e(al_b8da0e9e),
    .o(al_e94a3a72[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_76328905 (
    .a(al_9cdd3a01[0]),
    .b(al_9cdd3a01[1]),
    .c(al_9cdd3a01[2]),
    .d(al_9cdd3a01[3]),
    .e(al_9cdd3a01[4]),
    .f(al_b8da0e9e),
    .o(al_e94a3a72[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3bb7fc58 (
    .di(al_31a3e7af[125:124]),
    .raddr(al_e94a3a72),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_1591047a),
    .rdo(al_955db046[125:124]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d2f8de91 (
    .di(al_31a3e7af[123:122]),
    .raddr(al_e94a3a72),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_1591047a),
    .rdo(al_955db046[123:122]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_8c725d22 (
    .di(al_31a3e7af[121:120]),
    .raddr(al_e94a3a72),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_1591047a),
    .rdo(al_955db046[121:120]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_aa2c1e7 (
    .a(al_55ef04c8[0]),
    .b(al_fef4ecdb),
    .o(al_57782f22[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_938cc286 (
    .a(al_55ef04c8[0]),
    .b(al_55ef04c8[1]),
    .c(al_fef4ecdb),
    .o(al_57782f22[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_4745e6d3 (
    .a(al_55ef04c8[0]),
    .b(al_55ef04c8[1]),
    .c(al_55ef04c8[2]),
    .d(al_fef4ecdb),
    .o(al_57782f22[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_51aae568 (
    .a(al_55ef04c8[0]),
    .b(al_55ef04c8[1]),
    .c(al_55ef04c8[2]),
    .d(al_55ef04c8[3]),
    .e(al_fef4ecdb),
    .o(al_57782f22[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_aee99ad (
    .a(al_55ef04c8[0]),
    .b(al_55ef04c8[1]),
    .c(al_55ef04c8[2]),
    .d(al_55ef04c8[3]),
    .e(al_55ef04c8[4]),
    .f(al_fef4ecdb),
    .o(al_57782f22[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bb77db3f (
    .di(al_31a3e7af[131:130]),
    .raddr(al_57782f22),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d3c4d360),
    .rdo(al_955db046[131:130]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7a2809b8 (
    .di(al_31a3e7af[129:128]),
    .raddr(al_57782f22),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d3c4d360),
    .rdo(al_955db046[129:128]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e5bddef6 (
    .di(al_31a3e7af[127:126]),
    .raddr(al_57782f22),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d3c4d360),
    .rdo(al_955db046[127:126]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_deabc205 (
    .a(al_384dd51d[0]),
    .b(al_796e34c4),
    .o(al_9f1bb485[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_54995790 (
    .a(al_384dd51d[0]),
    .b(al_384dd51d[1]),
    .c(al_796e34c4),
    .o(al_9f1bb485[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_c396b12d (
    .a(al_384dd51d[0]),
    .b(al_384dd51d[1]),
    .c(al_384dd51d[2]),
    .d(al_796e34c4),
    .o(al_9f1bb485[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_beaa64c7 (
    .a(al_384dd51d[0]),
    .b(al_384dd51d[1]),
    .c(al_384dd51d[2]),
    .d(al_384dd51d[3]),
    .e(al_796e34c4),
    .o(al_9f1bb485[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_2545c3dd (
    .a(al_384dd51d[0]),
    .b(al_384dd51d[1]),
    .c(al_384dd51d[2]),
    .d(al_384dd51d[3]),
    .e(al_384dd51d[4]),
    .f(al_796e34c4),
    .o(al_9f1bb485[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e19f15ea (
    .di(al_31a3e7af[137:136]),
    .raddr(al_9f1bb485),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6d6760dd),
    .rdo(al_955db046[137:136]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e1f6a9f4 (
    .di(al_31a3e7af[135:134]),
    .raddr(al_9f1bb485),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6d6760dd),
    .rdo(al_955db046[135:134]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_91b97af1 (
    .di(al_31a3e7af[133:132]),
    .raddr(al_9f1bb485),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6d6760dd),
    .rdo(al_955db046[133:132]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_62e9c97d (
    .a(al_269b6545[0]),
    .b(al_df7aa915),
    .o(al_52fa7a1e[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_56a72c5e (
    .a(al_269b6545[0]),
    .b(al_269b6545[1]),
    .c(al_df7aa915),
    .o(al_52fa7a1e[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_7a132259 (
    .a(al_269b6545[0]),
    .b(al_269b6545[1]),
    .c(al_269b6545[2]),
    .d(al_df7aa915),
    .o(al_52fa7a1e[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_7e3a018b (
    .a(al_269b6545[0]),
    .b(al_269b6545[1]),
    .c(al_269b6545[2]),
    .d(al_269b6545[3]),
    .e(al_df7aa915),
    .o(al_52fa7a1e[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_bd7447f7 (
    .a(al_269b6545[0]),
    .b(al_269b6545[1]),
    .c(al_269b6545[2]),
    .d(al_269b6545[3]),
    .e(al_269b6545[4]),
    .f(al_df7aa915),
    .o(al_52fa7a1e[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f99bce81 (
    .di(al_31a3e7af[143:142]),
    .raddr(al_52fa7a1e),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_9cf6a965),
    .rdo(al_955db046[143:142]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7bb620ec (
    .di(al_31a3e7af[141:140]),
    .raddr(al_52fa7a1e),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_9cf6a965),
    .rdo(al_955db046[141:140]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_6477a992 (
    .di(al_31a3e7af[139:138]),
    .raddr(al_52fa7a1e),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_9cf6a965),
    .rdo(al_955db046[139:138]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_16f07168 (
    .a(al_430dd919[0]),
    .b(al_6dc98a03),
    .o(al_b81cf447[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_1314c625 (
    .a(al_430dd919[0]),
    .b(al_430dd919[1]),
    .c(al_6dc98a03),
    .o(al_b81cf447[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_4804d752 (
    .a(al_430dd919[0]),
    .b(al_430dd919[1]),
    .c(al_430dd919[2]),
    .d(al_6dc98a03),
    .o(al_b81cf447[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_47439294 (
    .a(al_430dd919[0]),
    .b(al_430dd919[1]),
    .c(al_430dd919[2]),
    .d(al_430dd919[3]),
    .e(al_6dc98a03),
    .o(al_b81cf447[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_edb17f8d (
    .a(al_430dd919[0]),
    .b(al_430dd919[1]),
    .c(al_430dd919[2]),
    .d(al_430dd919[3]),
    .e(al_430dd919[4]),
    .f(al_6dc98a03),
    .o(al_b81cf447[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_805fdbac (
    .di(al_31a3e7af[149:148]),
    .raddr(al_b81cf447),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_37a8c4a3),
    .rdo(al_955db046[149:148]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_af5fb389 (
    .di(al_31a3e7af[147:146]),
    .raddr(al_b81cf447),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_37a8c4a3),
    .rdo(al_955db046[147:146]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_464458d5 (
    .di(al_31a3e7af[145:144]),
    .raddr(al_b81cf447),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_37a8c4a3),
    .rdo(al_955db046[145:144]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_796ac887 (
    .a(al_5c6ba19f[0]),
    .b(al_80360204),
    .o(al_5fdc2ca7[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_a90fb196 (
    .a(al_5c6ba19f[0]),
    .b(al_5c6ba19f[1]),
    .c(al_80360204),
    .o(al_5fdc2ca7[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_3a9f58a9 (
    .a(al_5c6ba19f[0]),
    .b(al_5c6ba19f[1]),
    .c(al_5c6ba19f[2]),
    .d(al_80360204),
    .o(al_5fdc2ca7[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_cccf8488 (
    .a(al_5c6ba19f[0]),
    .b(al_5c6ba19f[1]),
    .c(al_5c6ba19f[2]),
    .d(al_5c6ba19f[3]),
    .e(al_80360204),
    .o(al_5fdc2ca7[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_747dc0b4 (
    .a(al_5c6ba19f[0]),
    .b(al_5c6ba19f[1]),
    .c(al_5c6ba19f[2]),
    .d(al_5c6ba19f[3]),
    .e(al_5c6ba19f[4]),
    .f(al_80360204),
    .o(al_5fdc2ca7[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_8b4a5b7f (
    .di(al_31a3e7af[155:154]),
    .raddr(al_5fdc2ca7),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2c31bcd7),
    .rdo(al_955db046[155:154]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b541b966 (
    .di(al_31a3e7af[153:152]),
    .raddr(al_5fdc2ca7),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2c31bcd7),
    .rdo(al_955db046[153:152]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bb14afba (
    .di(al_31a3e7af[151:150]),
    .raddr(al_5fdc2ca7),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2c31bcd7),
    .rdo(al_955db046[151:150]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_24406f19 (
    .a(al_4f6bae56[0]),
    .b(al_2bb74c3d),
    .o(al_2ad878de[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_a726b5a7 (
    .a(al_4f6bae56[0]),
    .b(al_4f6bae56[1]),
    .c(al_2bb74c3d),
    .o(al_2ad878de[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_f28ad40 (
    .a(al_4f6bae56[0]),
    .b(al_4f6bae56[1]),
    .c(al_4f6bae56[2]),
    .d(al_2bb74c3d),
    .o(al_2ad878de[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_46cb6c24 (
    .a(al_4f6bae56[0]),
    .b(al_4f6bae56[1]),
    .c(al_4f6bae56[2]),
    .d(al_4f6bae56[3]),
    .e(al_2bb74c3d),
    .o(al_2ad878de[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_528bca39 (
    .a(al_4f6bae56[0]),
    .b(al_4f6bae56[1]),
    .c(al_4f6bae56[2]),
    .d(al_4f6bae56[3]),
    .e(al_4f6bae56[4]),
    .f(al_2bb74c3d),
    .o(al_2ad878de[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_5c9c3cc7 (
    .di(al_31a3e7af[161:160]),
    .raddr(al_2ad878de),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_bbe31482),
    .rdo(al_955db046[161:160]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c4776815 (
    .di(al_31a3e7af[159:158]),
    .raddr(al_2ad878de),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_bbe31482),
    .rdo(al_955db046[159:158]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d5a897c2 (
    .di(al_31a3e7af[157:156]),
    .raddr(al_2ad878de),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_bbe31482),
    .rdo(al_955db046[157:156]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_7fdd4419 (
    .a(al_206e4ef2[0]),
    .b(al_9dcab982),
    .o(al_9ef91e29[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_33c2c060 (
    .a(al_206e4ef2[0]),
    .b(al_206e4ef2[1]),
    .c(al_9dcab982),
    .o(al_9ef91e29[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_225b14aa (
    .a(al_206e4ef2[0]),
    .b(al_206e4ef2[1]),
    .c(al_206e4ef2[2]),
    .d(al_9dcab982),
    .o(al_9ef91e29[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_73f895fa (
    .a(al_206e4ef2[0]),
    .b(al_206e4ef2[1]),
    .c(al_206e4ef2[2]),
    .d(al_206e4ef2[3]),
    .e(al_9dcab982),
    .o(al_9ef91e29[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_e1d44ab5 (
    .a(al_206e4ef2[0]),
    .b(al_206e4ef2[1]),
    .c(al_206e4ef2[2]),
    .d(al_206e4ef2[3]),
    .e(al_206e4ef2[4]),
    .f(al_9dcab982),
    .o(al_9ef91e29[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7fe34f12 (
    .di(al_31a3e7af[167:166]),
    .raddr(al_9ef91e29),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_edff11e6),
    .rdo(al_955db046[167:166]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_4d0f065d (
    .di(al_31a3e7af[165:164]),
    .raddr(al_9ef91e29),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_edff11e6),
    .rdo(al_955db046[165:164]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_10875757 (
    .di(al_31a3e7af[163:162]),
    .raddr(al_9ef91e29),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_edff11e6),
    .rdo(al_955db046[163:162]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_230ce711 (
    .a(al_ead25ba5[0]),
    .b(al_a9490be8),
    .o(al_b1ca7bde[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_ff1f4c3f (
    .a(al_ead25ba5[0]),
    .b(al_ead25ba5[1]),
    .c(al_a9490be8),
    .o(al_b1ca7bde[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_a6689926 (
    .a(al_ead25ba5[0]),
    .b(al_ead25ba5[1]),
    .c(al_ead25ba5[2]),
    .d(al_a9490be8),
    .o(al_b1ca7bde[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_226ccfb5 (
    .a(al_ead25ba5[0]),
    .b(al_ead25ba5[1]),
    .c(al_ead25ba5[2]),
    .d(al_ead25ba5[3]),
    .e(al_a9490be8),
    .o(al_b1ca7bde[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_aa5d5ec3 (
    .a(al_ead25ba5[0]),
    .b(al_ead25ba5[1]),
    .c(al_ead25ba5[2]),
    .d(al_ead25ba5[3]),
    .e(al_ead25ba5[4]),
    .f(al_a9490be8),
    .o(al_b1ca7bde[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b90b2c0b (
    .di(al_31a3e7af[173:172]),
    .raddr(al_b1ca7bde),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_4b287773),
    .rdo(al_955db046[173:172]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_375ec505 (
    .di(al_31a3e7af[171:170]),
    .raddr(al_b1ca7bde),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_4b287773),
    .rdo(al_955db046[171:170]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_727c3adb (
    .di(al_31a3e7af[169:168]),
    .raddr(al_b1ca7bde),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_4b287773),
    .rdo(al_955db046[169:168]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_6acf04a5 (
    .a(al_b04a4cbc[0]),
    .b(al_28d8d34d),
    .o(al_54ef982d[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_bfd63925 (
    .a(al_b04a4cbc[0]),
    .b(al_b04a4cbc[1]),
    .c(al_28d8d34d),
    .o(al_54ef982d[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_bf19a826 (
    .a(al_b04a4cbc[0]),
    .b(al_b04a4cbc[1]),
    .c(al_b04a4cbc[2]),
    .d(al_28d8d34d),
    .o(al_54ef982d[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_917c7de3 (
    .a(al_b04a4cbc[0]),
    .b(al_b04a4cbc[1]),
    .c(al_b04a4cbc[2]),
    .d(al_b04a4cbc[3]),
    .e(al_28d8d34d),
    .o(al_54ef982d[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_c5f5c704 (
    .a(al_b04a4cbc[0]),
    .b(al_b04a4cbc[1]),
    .c(al_b04a4cbc[2]),
    .d(al_b04a4cbc[3]),
    .e(al_b04a4cbc[4]),
    .f(al_28d8d34d),
    .o(al_54ef982d[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c73033c4 (
    .di(al_31a3e7af[179:178]),
    .raddr(al_54ef982d),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_a18a78ec),
    .rdo(al_955db046[179:178]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9e9eaefb (
    .di(al_31a3e7af[177:176]),
    .raddr(al_54ef982d),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_a18a78ec),
    .rdo(al_955db046[177:176]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_6ef12f18 (
    .di(al_31a3e7af[175:174]),
    .raddr(al_54ef982d),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_a18a78ec),
    .rdo(al_955db046[175:174]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_486f21c5 (
    .a(al_6b9e1d84[0]),
    .b(al_e6ea44e6),
    .o(al_84ba38ec[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_9403205f (
    .a(al_6b9e1d84[0]),
    .b(al_6b9e1d84[1]),
    .c(al_e6ea44e6),
    .o(al_84ba38ec[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_f7d1a670 (
    .a(al_6b9e1d84[0]),
    .b(al_6b9e1d84[1]),
    .c(al_6b9e1d84[2]),
    .d(al_e6ea44e6),
    .o(al_84ba38ec[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_da642c00 (
    .a(al_6b9e1d84[0]),
    .b(al_6b9e1d84[1]),
    .c(al_6b9e1d84[2]),
    .d(al_6b9e1d84[3]),
    .e(al_e6ea44e6),
    .o(al_84ba38ec[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_1b480f6e (
    .a(al_6b9e1d84[0]),
    .b(al_6b9e1d84[1]),
    .c(al_6b9e1d84[2]),
    .d(al_6b9e1d84[3]),
    .e(al_6b9e1d84[4]),
    .f(al_e6ea44e6),
    .o(al_84ba38ec[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_53910f01 (
    .di(al_31a3e7af[17:16]),
    .raddr(al_84ba38ec),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f8b11b95),
    .rdo(al_955db046[17:16]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_4178ae2f (
    .di(al_31a3e7af[15:14]),
    .raddr(al_84ba38ec),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f8b11b95),
    .rdo(al_955db046[15:14]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_4c21553b (
    .di(al_31a3e7af[13:12]),
    .raddr(al_84ba38ec),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f8b11b95),
    .rdo(al_955db046[13:12]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_eca00686 (
    .a(al_c244bf8b[0]),
    .b(al_7cd149c6),
    .o(al_8bf0a0c9[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_422adb3f (
    .a(al_c244bf8b[0]),
    .b(al_c244bf8b[1]),
    .c(al_7cd149c6),
    .o(al_8bf0a0c9[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_b9531746 (
    .a(al_c244bf8b[0]),
    .b(al_c244bf8b[1]),
    .c(al_c244bf8b[2]),
    .d(al_7cd149c6),
    .o(al_8bf0a0c9[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_400e74f5 (
    .a(al_c244bf8b[0]),
    .b(al_c244bf8b[1]),
    .c(al_c244bf8b[2]),
    .d(al_c244bf8b[3]),
    .e(al_7cd149c6),
    .o(al_8bf0a0c9[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_a7bf22f (
    .a(al_c244bf8b[0]),
    .b(al_c244bf8b[1]),
    .c(al_c244bf8b[2]),
    .d(al_c244bf8b[3]),
    .e(al_c244bf8b[4]),
    .f(al_7cd149c6),
    .o(al_8bf0a0c9[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_25cdd519 (
    .di(al_31a3e7af[185:184]),
    .raddr(al_8bf0a0c9),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_dd0c66b3),
    .rdo(al_955db046[185:184]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_96bed03a (
    .di(al_31a3e7af[183:182]),
    .raddr(al_8bf0a0c9),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_dd0c66b3),
    .rdo(al_955db046[183:182]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_30ef8598 (
    .di(al_31a3e7af[181:180]),
    .raddr(al_8bf0a0c9),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_dd0c66b3),
    .rdo(al_955db046[181:180]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_71bf9757 (
    .a(al_d44a73a0[0]),
    .b(al_b56307ec),
    .o(al_cb2afcca[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_32cd6c01 (
    .a(al_d44a73a0[0]),
    .b(al_d44a73a0[1]),
    .c(al_b56307ec),
    .o(al_cb2afcca[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_811b1668 (
    .a(al_d44a73a0[0]),
    .b(al_d44a73a0[1]),
    .c(al_d44a73a0[2]),
    .d(al_b56307ec),
    .o(al_cb2afcca[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_67cf69f0 (
    .a(al_d44a73a0[0]),
    .b(al_d44a73a0[1]),
    .c(al_d44a73a0[2]),
    .d(al_d44a73a0[3]),
    .e(al_b56307ec),
    .o(al_cb2afcca[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_b0b3c5ec (
    .a(al_d44a73a0[0]),
    .b(al_d44a73a0[1]),
    .c(al_d44a73a0[2]),
    .d(al_d44a73a0[3]),
    .e(al_d44a73a0[4]),
    .f(al_b56307ec),
    .o(al_cb2afcca[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9811c5a (
    .di(al_31a3e7af[191:190]),
    .raddr(al_cb2afcca),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_edb83574),
    .rdo(al_955db046[191:190]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_16c38ff3 (
    .di(al_31a3e7af[189:188]),
    .raddr(al_cb2afcca),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_edb83574),
    .rdo(al_955db046[189:188]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_627b8304 (
    .di(al_31a3e7af[187:186]),
    .raddr(al_cb2afcca),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_edb83574),
    .rdo(al_955db046[187:186]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_5889d043 (
    .a(al_37663fe4[0]),
    .b(al_31be1d74),
    .o(al_43333b4e[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_89d38d89 (
    .a(al_37663fe4[0]),
    .b(al_37663fe4[1]),
    .c(al_31be1d74),
    .o(al_43333b4e[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_c2154b65 (
    .a(al_37663fe4[0]),
    .b(al_37663fe4[1]),
    .c(al_37663fe4[2]),
    .d(al_31be1d74),
    .o(al_43333b4e[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_74152eaf (
    .a(al_37663fe4[0]),
    .b(al_37663fe4[1]),
    .c(al_37663fe4[2]),
    .d(al_37663fe4[3]),
    .e(al_31be1d74),
    .o(al_43333b4e[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_a8cc5672 (
    .a(al_37663fe4[0]),
    .b(al_37663fe4[1]),
    .c(al_37663fe4[2]),
    .d(al_37663fe4[3]),
    .e(al_37663fe4[4]),
    .f(al_31be1d74),
    .o(al_43333b4e[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_208e4cfe (
    .di(al_31a3e7af[197:196]),
    .raddr(al_43333b4e),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2935d0ed),
    .rdo(al_955db046[197:196]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_6b691fc1 (
    .di(al_31a3e7af[195:194]),
    .raddr(al_43333b4e),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2935d0ed),
    .rdo(al_955db046[195:194]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3e62c713 (
    .di(al_31a3e7af[193:192]),
    .raddr(al_43333b4e),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2935d0ed),
    .rdo(al_955db046[193:192]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_808e6380 (
    .a(al_e865b87a[0]),
    .b(al_cc2e5bcc),
    .o(al_ad11f805[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_3d300dee (
    .a(al_e865b87a[0]),
    .b(al_e865b87a[1]),
    .c(al_cc2e5bcc),
    .o(al_ad11f805[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_c2a1213f (
    .a(al_e865b87a[0]),
    .b(al_e865b87a[1]),
    .c(al_e865b87a[2]),
    .d(al_cc2e5bcc),
    .o(al_ad11f805[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_210e3038 (
    .a(al_e865b87a[0]),
    .b(al_e865b87a[1]),
    .c(al_e865b87a[2]),
    .d(al_e865b87a[3]),
    .e(al_cc2e5bcc),
    .o(al_ad11f805[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_52ba792b (
    .a(al_e865b87a[0]),
    .b(al_e865b87a[1]),
    .c(al_e865b87a[2]),
    .d(al_e865b87a[3]),
    .e(al_e865b87a[4]),
    .f(al_cc2e5bcc),
    .o(al_ad11f805[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c788c834 (
    .di(al_31a3e7af[203:202]),
    .raddr(al_ad11f805),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_538eda90),
    .rdo(al_955db046[203:202]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bc4763b7 (
    .di(al_31a3e7af[201:200]),
    .raddr(al_ad11f805),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_538eda90),
    .rdo(al_955db046[201:200]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7a9a445b (
    .di(al_31a3e7af[199:198]),
    .raddr(al_ad11f805),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_538eda90),
    .rdo(al_955db046[199:198]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_357d3c57 (
    .a(al_f359f0c8[0]),
    .b(al_ee615f87),
    .o(al_e4f3a09c[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_a5e60d7f (
    .a(al_f359f0c8[0]),
    .b(al_f359f0c8[1]),
    .c(al_ee615f87),
    .o(al_e4f3a09c[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_30bf13dc (
    .a(al_f359f0c8[0]),
    .b(al_f359f0c8[1]),
    .c(al_f359f0c8[2]),
    .d(al_ee615f87),
    .o(al_e4f3a09c[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_f2bfb6e3 (
    .a(al_f359f0c8[0]),
    .b(al_f359f0c8[1]),
    .c(al_f359f0c8[2]),
    .d(al_f359f0c8[3]),
    .e(al_ee615f87),
    .o(al_e4f3a09c[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_81816f43 (
    .a(al_f359f0c8[0]),
    .b(al_f359f0c8[1]),
    .c(al_f359f0c8[2]),
    .d(al_f359f0c8[3]),
    .e(al_f359f0c8[4]),
    .f(al_ee615f87),
    .o(al_e4f3a09c[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ea6d15af (
    .di(al_31a3e7af[209:208]),
    .raddr(al_e4f3a09c),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2503fdb),
    .rdo(al_955db046[209:208]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d4e09a27 (
    .di(al_31a3e7af[207:206]),
    .raddr(al_e4f3a09c),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2503fdb),
    .rdo(al_955db046[207:206]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_31f9dc84 (
    .di(al_31a3e7af[205:204]),
    .raddr(al_e4f3a09c),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_2503fdb),
    .rdo(al_955db046[205:204]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_bfac78ce (
    .a(al_85a14e36[0]),
    .b(al_35f768f4),
    .o(al_eb6aa70a[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_d3e662db (
    .a(al_85a14e36[0]),
    .b(al_85a14e36[1]),
    .c(al_35f768f4),
    .o(al_eb6aa70a[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_db541318 (
    .a(al_85a14e36[0]),
    .b(al_85a14e36[1]),
    .c(al_85a14e36[2]),
    .d(al_35f768f4),
    .o(al_eb6aa70a[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_35ffa9a1 (
    .a(al_85a14e36[0]),
    .b(al_85a14e36[1]),
    .c(al_85a14e36[2]),
    .d(al_85a14e36[3]),
    .e(al_35f768f4),
    .o(al_eb6aa70a[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_cbd0b568 (
    .a(al_85a14e36[0]),
    .b(al_85a14e36[1]),
    .c(al_85a14e36[2]),
    .d(al_85a14e36[3]),
    .e(al_85a14e36[4]),
    .f(al_35f768f4),
    .o(al_eb6aa70a[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ef1df979 (
    .di(al_31a3e7af[215:214]),
    .raddr(al_eb6aa70a),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f8fcd204),
    .rdo(al_955db046[215:214]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bccd32bb (
    .di(al_31a3e7af[213:212]),
    .raddr(al_eb6aa70a),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f8fcd204),
    .rdo(al_955db046[213:212]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c580087a (
    .di(al_31a3e7af[211:210]),
    .raddr(al_eb6aa70a),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f8fcd204),
    .rdo(al_955db046[211:210]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_b32d4cf2 (
    .a(al_e31889d8[0]),
    .b(al_5e6f3859),
    .o(al_6101d7c8[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_93009c2e (
    .a(al_e31889d8[0]),
    .b(al_e31889d8[1]),
    .c(al_5e6f3859),
    .o(al_6101d7c8[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_347dab58 (
    .a(al_e31889d8[0]),
    .b(al_e31889d8[1]),
    .c(al_e31889d8[2]),
    .d(al_5e6f3859),
    .o(al_6101d7c8[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_eb62178 (
    .a(al_e31889d8[0]),
    .b(al_e31889d8[1]),
    .c(al_e31889d8[2]),
    .d(al_e31889d8[3]),
    .e(al_5e6f3859),
    .o(al_6101d7c8[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_2329bc9e (
    .a(al_e31889d8[0]),
    .b(al_e31889d8[1]),
    .c(al_e31889d8[2]),
    .d(al_e31889d8[3]),
    .e(al_e31889d8[4]),
    .f(al_5e6f3859),
    .o(al_6101d7c8[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_6784ac34 (
    .di(al_31a3e7af[221:220]),
    .raddr(al_6101d7c8),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_467a2ca),
    .rdo(al_955db046[221:220]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_dcb19d9e (
    .di(al_31a3e7af[219:218]),
    .raddr(al_6101d7c8),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_467a2ca),
    .rdo(al_955db046[219:218]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2f5250f4 (
    .di(al_31a3e7af[217:216]),
    .raddr(al_6101d7c8),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_467a2ca),
    .rdo(al_955db046[217:216]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_31e2b01c (
    .a(al_8349e0d1[0]),
    .b(al_2efa36ca),
    .o(al_9bd5fcab[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_274609c5 (
    .a(al_8349e0d1[0]),
    .b(al_8349e0d1[1]),
    .c(al_2efa36ca),
    .o(al_9bd5fcab[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_6a06b423 (
    .a(al_8349e0d1[0]),
    .b(al_8349e0d1[1]),
    .c(al_8349e0d1[2]),
    .d(al_2efa36ca),
    .o(al_9bd5fcab[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_790665d9 (
    .a(al_8349e0d1[0]),
    .b(al_8349e0d1[1]),
    .c(al_8349e0d1[2]),
    .d(al_8349e0d1[3]),
    .e(al_2efa36ca),
    .o(al_9bd5fcab[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_403cce4c (
    .a(al_8349e0d1[0]),
    .b(al_8349e0d1[1]),
    .c(al_8349e0d1[2]),
    .d(al_8349e0d1[3]),
    .e(al_8349e0d1[4]),
    .f(al_2efa36ca),
    .o(al_9bd5fcab[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c1d26866 (
    .di(al_31a3e7af[227:226]),
    .raddr(al_9bd5fcab),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_c76ae5c3),
    .rdo(al_955db046[227:226]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_72a3c983 (
    .di(al_31a3e7af[225:224]),
    .raddr(al_9bd5fcab),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_c76ae5c3),
    .rdo(al_955db046[225:224]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_fc65d58f (
    .di(al_31a3e7af[223:222]),
    .raddr(al_9bd5fcab),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_c76ae5c3),
    .rdo(al_955db046[223:222]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_32bbfc5b (
    .a(al_2ef171e7[0]),
    .b(al_4708b339),
    .o(al_c408b364[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_f104a34a (
    .a(al_2ef171e7[0]),
    .b(al_2ef171e7[1]),
    .c(al_4708b339),
    .o(al_c408b364[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_83c13b02 (
    .a(al_2ef171e7[0]),
    .b(al_2ef171e7[1]),
    .c(al_2ef171e7[2]),
    .d(al_4708b339),
    .o(al_c408b364[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_2d9a943d (
    .a(al_2ef171e7[0]),
    .b(al_2ef171e7[1]),
    .c(al_2ef171e7[2]),
    .d(al_2ef171e7[3]),
    .e(al_4708b339),
    .o(al_c408b364[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_f150976e (
    .a(al_2ef171e7[0]),
    .b(al_2ef171e7[1]),
    .c(al_2ef171e7[2]),
    .d(al_2ef171e7[3]),
    .e(al_2ef171e7[4]),
    .f(al_4708b339),
    .o(al_c408b364[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_70d1724c (
    .di(al_31a3e7af[233:232]),
    .raddr(al_c408b364),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d2c8f1b1),
    .rdo(al_955db046[233:232]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_92709234 (
    .di(al_31a3e7af[231:230]),
    .raddr(al_c408b364),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d2c8f1b1),
    .rdo(al_955db046[231:230]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bad7713d (
    .di(al_31a3e7af[229:228]),
    .raddr(al_c408b364),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d2c8f1b1),
    .rdo(al_955db046[229:228]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_bb22d794 (
    .a(al_662b3089[0]),
    .b(al_4864d933),
    .o(al_b96545cc[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_21913106 (
    .a(al_662b3089[0]),
    .b(al_662b3089[1]),
    .c(al_4864d933),
    .o(al_b96545cc[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_7406ba (
    .a(al_662b3089[0]),
    .b(al_662b3089[1]),
    .c(al_662b3089[2]),
    .d(al_4864d933),
    .o(al_b96545cc[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_3f4d90ce (
    .a(al_662b3089[0]),
    .b(al_662b3089[1]),
    .c(al_662b3089[2]),
    .d(al_662b3089[3]),
    .e(al_4864d933),
    .o(al_b96545cc[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_5e0b0e75 (
    .a(al_662b3089[0]),
    .b(al_662b3089[1]),
    .c(al_662b3089[2]),
    .d(al_662b3089[3]),
    .e(al_662b3089[4]),
    .f(al_4864d933),
    .o(al_b96545cc[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_360d52fe (
    .di(al_31a3e7af[239:238]),
    .raddr(al_b96545cc),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_282d371d),
    .rdo(al_955db046[239:238]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_eccca561 (
    .di(al_31a3e7af[237:236]),
    .raddr(al_b96545cc),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_282d371d),
    .rdo(al_955db046[237:236]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2a22c18d (
    .di(al_31a3e7af[235:234]),
    .raddr(al_b96545cc),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_282d371d),
    .rdo(al_955db046[235:234]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_bb93b4a3 (
    .a(al_4a30bd0f[0]),
    .b(al_71cac35e),
    .o(al_556b029f[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_e54050ea (
    .a(al_4a30bd0f[0]),
    .b(al_4a30bd0f[1]),
    .c(al_71cac35e),
    .o(al_556b029f[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_62880ef3 (
    .a(al_4a30bd0f[0]),
    .b(al_4a30bd0f[1]),
    .c(al_4a30bd0f[2]),
    .d(al_71cac35e),
    .o(al_556b029f[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_d32fe990 (
    .a(al_4a30bd0f[0]),
    .b(al_4a30bd0f[1]),
    .c(al_4a30bd0f[2]),
    .d(al_4a30bd0f[3]),
    .e(al_71cac35e),
    .o(al_556b029f[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_c7d24859 (
    .a(al_4a30bd0f[0]),
    .b(al_4a30bd0f[1]),
    .c(al_4a30bd0f[2]),
    .d(al_4a30bd0f[3]),
    .e(al_4a30bd0f[4]),
    .f(al_71cac35e),
    .o(al_556b029f[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9d5f12f5 (
    .di(al_31a3e7af[23:22]),
    .raddr(al_556b029f),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_cd27f05c),
    .rdo(al_955db046[23:22]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_64bcb047 (
    .di(al_31a3e7af[21:20]),
    .raddr(al_556b029f),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_cd27f05c),
    .rdo(al_955db046[21:20]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_8dc13ea4 (
    .di(al_31a3e7af[19:18]),
    .raddr(al_556b029f),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_cd27f05c),
    .rdo(al_955db046[19:18]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_8ad037ce (
    .a(al_2119f32d[0]),
    .b(al_c3e70575),
    .o(al_4f1aa340[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_40e8a54c (
    .a(al_2119f32d[0]),
    .b(al_2119f32d[1]),
    .c(al_c3e70575),
    .o(al_4f1aa340[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_d86f4356 (
    .a(al_2119f32d[0]),
    .b(al_2119f32d[1]),
    .c(al_2119f32d[2]),
    .d(al_c3e70575),
    .o(al_4f1aa340[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_8e6069b4 (
    .a(al_2119f32d[0]),
    .b(al_2119f32d[1]),
    .c(al_2119f32d[2]),
    .d(al_2119f32d[3]),
    .e(al_c3e70575),
    .o(al_4f1aa340[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_733985d0 (
    .a(al_2119f32d[0]),
    .b(al_2119f32d[1]),
    .c(al_2119f32d[2]),
    .d(al_2119f32d[3]),
    .e(al_2119f32d[4]),
    .f(al_c3e70575),
    .o(al_4f1aa340[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_19a1fe7a (
    .di(al_31a3e7af[245:244]),
    .raddr(al_4f1aa340),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_27b77d58),
    .rdo(al_955db046[245:244]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_92b3968e (
    .di(al_31a3e7af[243:242]),
    .raddr(al_4f1aa340),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_27b77d58),
    .rdo(al_955db046[243:242]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_fbf6fbef (
    .di(al_31a3e7af[241:240]),
    .raddr(al_4f1aa340),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_27b77d58),
    .rdo(al_955db046[241:240]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e83aedd4 (
    .a(al_d9591ec3[0]),
    .b(al_83ebd977),
    .o(al_902090d1[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_f823ec51 (
    .a(al_d9591ec3[0]),
    .b(al_d9591ec3[1]),
    .c(al_83ebd977),
    .o(al_902090d1[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_f34148ba (
    .a(al_d9591ec3[0]),
    .b(al_d9591ec3[1]),
    .c(al_d9591ec3[2]),
    .d(al_83ebd977),
    .o(al_902090d1[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_b1f44fa6 (
    .a(al_d9591ec3[0]),
    .b(al_d9591ec3[1]),
    .c(al_d9591ec3[2]),
    .d(al_d9591ec3[3]),
    .e(al_83ebd977),
    .o(al_902090d1[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_2826a8b8 (
    .a(al_d9591ec3[0]),
    .b(al_d9591ec3[1]),
    .c(al_d9591ec3[2]),
    .d(al_d9591ec3[3]),
    .e(al_d9591ec3[4]),
    .f(al_83ebd977),
    .o(al_902090d1[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_8330c5d7 (
    .di(al_31a3e7af[251:250]),
    .raddr(al_902090d1),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d4d145cc),
    .rdo(al_955db046[251:250]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c5b91ab7 (
    .di(al_31a3e7af[249:248]),
    .raddr(al_902090d1),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d4d145cc),
    .rdo(al_955db046[249:248]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_aa4a6cce (
    .di(al_31a3e7af[247:246]),
    .raddr(al_902090d1),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_d4d145cc),
    .rdo(al_955db046[247:246]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_5c3d1d4a (
    .a(al_1d102248[0]),
    .b(al_6bddd01a),
    .o(al_2e33811d[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_f962ad77 (
    .a(al_1d102248[0]),
    .b(al_1d102248[1]),
    .c(al_6bddd01a),
    .o(al_2e33811d[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_130218c3 (
    .a(al_1d102248[0]),
    .b(al_1d102248[1]),
    .c(al_1d102248[2]),
    .d(al_6bddd01a),
    .o(al_2e33811d[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_a995f945 (
    .a(al_1d102248[0]),
    .b(al_1d102248[1]),
    .c(al_1d102248[2]),
    .d(al_1d102248[3]),
    .e(al_6bddd01a),
    .o(al_2e33811d[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_da0a03db (
    .a(al_1d102248[0]),
    .b(al_1d102248[1]),
    .c(al_1d102248[2]),
    .d(al_1d102248[3]),
    .e(al_1d102248[4]),
    .f(al_6bddd01a),
    .o(al_2e33811d[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_6d1d7436 (
    .di(al_31a3e7af[255:254]),
    .raddr(al_2e33811d),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_129a2529),
    .rdo(al_955db046[255:254]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_db47d543 (
    .di(al_31a3e7af[253:252]),
    .raddr(al_2e33811d),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_129a2529),
    .rdo(al_955db046[253:252]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_5651af64 (
    .a(al_f78383db[0]),
    .b(al_c85cbcb),
    .o(al_6ab65bb5[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_7b1658c8 (
    .a(al_f78383db[0]),
    .b(al_f78383db[1]),
    .c(al_c85cbcb),
    .o(al_6ab65bb5[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_bbef904 (
    .a(al_f78383db[0]),
    .b(al_f78383db[1]),
    .c(al_f78383db[2]),
    .d(al_c85cbcb),
    .o(al_6ab65bb5[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_c3587a03 (
    .a(al_f78383db[0]),
    .b(al_f78383db[1]),
    .c(al_f78383db[2]),
    .d(al_f78383db[3]),
    .e(al_c85cbcb),
    .o(al_6ab65bb5[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_61fcd52d (
    .a(al_f78383db[0]),
    .b(al_f78383db[1]),
    .c(al_f78383db[2]),
    .d(al_f78383db[3]),
    .e(al_f78383db[4]),
    .f(al_c85cbcb),
    .o(al_6ab65bb5[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_45ccd5e1 (
    .di(al_31a3e7af[29:28]),
    .raddr(al_6ab65bb5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_14cefac2),
    .rdo(al_955db046[29:28]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_678d1b61 (
    .di(al_31a3e7af[27:26]),
    .raddr(al_6ab65bb5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_14cefac2),
    .rdo(al_955db046[27:26]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d4d7cb29 (
    .di(al_31a3e7af[25:24]),
    .raddr(al_6ab65bb5),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_14cefac2),
    .rdo(al_955db046[25:24]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_3446483 (
    .a(al_d9be1f39[0]),
    .b(al_f7c9608b),
    .o(al_8abfbd08[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_c301b328 (
    .a(al_d9be1f39[0]),
    .b(al_d9be1f39[1]),
    .c(al_f7c9608b),
    .o(al_8abfbd08[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_b3a182 (
    .a(al_d9be1f39[0]),
    .b(al_d9be1f39[1]),
    .c(al_d9be1f39[2]),
    .d(al_f7c9608b),
    .o(al_8abfbd08[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_634a9597 (
    .a(al_d9be1f39[0]),
    .b(al_d9be1f39[1]),
    .c(al_d9be1f39[2]),
    .d(al_d9be1f39[3]),
    .e(al_f7c9608b),
    .o(al_8abfbd08[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_b66d5934 (
    .a(al_d9be1f39[0]),
    .b(al_d9be1f39[1]),
    .c(al_d9be1f39[2]),
    .d(al_d9be1f39[3]),
    .e(al_d9be1f39[4]),
    .f(al_f7c9608b),
    .o(al_8abfbd08[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e71b06ef (
    .di(al_31a3e7af[35:34]),
    .raddr(al_8abfbd08),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6fd6ffff),
    .rdo(al_955db046[35:34]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_4d322413 (
    .di(al_31a3e7af[33:32]),
    .raddr(al_8abfbd08),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6fd6ffff),
    .rdo(al_955db046[33:32]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f2a19bd3 (
    .di(al_31a3e7af[31:30]),
    .raddr(al_8abfbd08),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_6fd6ffff),
    .rdo(al_955db046[31:30]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_877b4364 (
    .a(al_1e255230[0]),
    .b(al_ac593c94),
    .o(al_1a0d603f[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_55ace221 (
    .a(al_1e255230[0]),
    .b(al_1e255230[1]),
    .c(al_ac593c94),
    .o(al_1a0d603f[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_f9dbdc57 (
    .a(al_1e255230[0]),
    .b(al_1e255230[1]),
    .c(al_1e255230[2]),
    .d(al_ac593c94),
    .o(al_1a0d603f[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_56b9294 (
    .a(al_1e255230[0]),
    .b(al_1e255230[1]),
    .c(al_1e255230[2]),
    .d(al_1e255230[3]),
    .e(al_ac593c94),
    .o(al_1a0d603f[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_b4b93314 (
    .a(al_1e255230[0]),
    .b(al_1e255230[1]),
    .c(al_1e255230[2]),
    .d(al_1e255230[3]),
    .e(al_1e255230[4]),
    .f(al_ac593c94),
    .o(al_1a0d603f[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_78e6f247 (
    .di(al_31a3e7af[41:40]),
    .raddr(al_1a0d603f),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f645b571),
    .rdo(al_955db046[41:40]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7edf6059 (
    .di(al_31a3e7af[39:38]),
    .raddr(al_1a0d603f),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f645b571),
    .rdo(al_955db046[39:38]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_edf8d835 (
    .di(al_31a3e7af[37:36]),
    .raddr(al_1a0d603f),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_f645b571),
    .rdo(al_955db046[37:36]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_1a63c9a2 (
    .a(al_d61bccef[0]),
    .b(al_ad58fbc9),
    .o(al_8f8431f6[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_199db13a (
    .a(al_d61bccef[0]),
    .b(al_d61bccef[1]),
    .c(al_ad58fbc9),
    .o(al_8f8431f6[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_e71ae6b5 (
    .a(al_d61bccef[0]),
    .b(al_d61bccef[1]),
    .c(al_d61bccef[2]),
    .d(al_ad58fbc9),
    .o(al_8f8431f6[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_336022f9 (
    .a(al_d61bccef[0]),
    .b(al_d61bccef[1]),
    .c(al_d61bccef[2]),
    .d(al_d61bccef[3]),
    .e(al_ad58fbc9),
    .o(al_8f8431f6[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_e4af6562 (
    .a(al_d61bccef[0]),
    .b(al_d61bccef[1]),
    .c(al_d61bccef[2]),
    .d(al_d61bccef[3]),
    .e(al_d61bccef[4]),
    .f(al_ad58fbc9),
    .o(al_8f8431f6[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b259a8a0 (
    .di(al_31a3e7af[47:46]),
    .raddr(al_8f8431f6),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_3419432c),
    .rdo(al_955db046[47:46]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d37790c2 (
    .di(al_31a3e7af[45:44]),
    .raddr(al_8f8431f6),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_3419432c),
    .rdo(al_955db046[45:44]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_85310eaf (
    .di(al_31a3e7af[43:42]),
    .raddr(al_8f8431f6),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_3419432c),
    .rdo(al_955db046[43:42]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_f22850 (
    .a(al_46e8788c[0]),
    .b(al_3d66f550),
    .o(al_91916c28[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_c927d2bb (
    .a(al_46e8788c[0]),
    .b(al_46e8788c[1]),
    .c(al_3d66f550),
    .o(al_91916c28[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_eb7e19a1 (
    .a(al_46e8788c[0]),
    .b(al_46e8788c[1]),
    .c(al_46e8788c[2]),
    .d(al_3d66f550),
    .o(al_91916c28[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_747539db (
    .a(al_46e8788c[0]),
    .b(al_46e8788c[1]),
    .c(al_46e8788c[2]),
    .d(al_46e8788c[3]),
    .e(al_3d66f550),
    .o(al_91916c28[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_ab4f7613 (
    .a(al_46e8788c[0]),
    .b(al_46e8788c[1]),
    .c(al_46e8788c[2]),
    .d(al_46e8788c[3]),
    .e(al_46e8788c[4]),
    .f(al_3d66f550),
    .o(al_91916c28[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2ea7cf1c (
    .di(al_31a3e7af[53:52]),
    .raddr(al_91916c28),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_b9e4ee74),
    .rdo(al_955db046[53:52]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3ec98672 (
    .di(al_31a3e7af[51:50]),
    .raddr(al_91916c28),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_b9e4ee74),
    .rdo(al_955db046[51:50]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_aaeafe5b (
    .di(al_31a3e7af[49:48]),
    .raddr(al_91916c28),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_b9e4ee74),
    .rdo(al_955db046[49:48]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_af410a (
    .a(al_56e72bf4[0]),
    .b(al_12b38499),
    .o(al_27625f51[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_17f5c9b1 (
    .a(al_56e72bf4[0]),
    .b(al_56e72bf4[1]),
    .c(al_12b38499),
    .o(al_27625f51[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_8aa75dee (
    .a(al_56e72bf4[0]),
    .b(al_56e72bf4[1]),
    .c(al_56e72bf4[2]),
    .d(al_12b38499),
    .o(al_27625f51[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_94b7a3d7 (
    .a(al_56e72bf4[0]),
    .b(al_56e72bf4[1]),
    .c(al_56e72bf4[2]),
    .d(al_56e72bf4[3]),
    .e(al_12b38499),
    .o(al_27625f51[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_6231d4f7 (
    .a(al_56e72bf4[0]),
    .b(al_56e72bf4[1]),
    .c(al_56e72bf4[2]),
    .d(al_56e72bf4[3]),
    .e(al_56e72bf4[4]),
    .f(al_12b38499),
    .o(al_27625f51[4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_117e1a35 (
    .di(al_31a3e7af[59:58]),
    .raddr(al_27625f51),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_4b747cba),
    .rdo(al_955db046[59:58]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2e3ce087 (
    .di(al_31a3e7af[57:56]),
    .raddr(al_27625f51),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_4b747cba),
    .rdo(al_955db046[57:56]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e5ff4bda (
    .di(al_31a3e7af[55:54]),
    .raddr(al_27625f51),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_511af127),
    .wclk(al_ef3696df[0]),
    .we(al_4b747cba),
    .rdo(al_955db046[55:54]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ab7482db (
    .i(al_26a2c365),
    .o(al_a0e1d396[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_bee333e6 (
    .i(al_a0e1d396[0]),
    .o(al_4b4a698a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ce851c9 (
    .i(al_33cf56b3),
    .o(al_a0e1d396[10]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_86e995a8 (
    .i(al_a0e1d396[10]),
    .o(al_b8cc00cf));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_e0cbd333 (
    .i(al_39705b9f),
    .o(al_a0e1d396[11]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_dcbffbaa (
    .i(al_a0e1d396[11]),
    .o(al_106fddab));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b1c764c7 (
    .i(al_860bc871),
    .o(al_a0e1d396[12]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6abc4aa3 (
    .i(al_a0e1d396[12]),
    .o(al_82133c54));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1cc3c9b6 (
    .i(al_eda53b41),
    .o(al_a0e1d396[13]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1d8c6429 (
    .i(al_a0e1d396[13]),
    .o(al_9f6750b6));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_67f99eeb (
    .i(al_8695553e),
    .o(al_a0e1d396[14]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_16e2c7c9 (
    .i(al_a0e1d396[14]),
    .o(al_21d51e65));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f2487c2f (
    .i(al_646f260c),
    .o(al_a0e1d396[15]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_25a70cdc (
    .i(al_a0e1d396[15]),
    .o(al_3da9562a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_6ead66e3 (
    .i(al_2c63960b),
    .o(al_a0e1d396[16]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a1844748 (
    .i(al_a0e1d396[16]),
    .o(al_d9d76d0a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ca823f4f (
    .i(al_cea991a),
    .o(al_a0e1d396[17]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_63d17660 (
    .i(al_a0e1d396[17]),
    .o(al_64f79045));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b616339 (
    .i(al_fdd1bba3),
    .o(al_a0e1d396[18]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1dd47a4a (
    .i(al_a0e1d396[18]),
    .o(al_ab1b2b16));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_fddad69 (
    .i(al_7ceaf80e),
    .o(al_a0e1d396[19]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2e89c5ef (
    .i(al_a0e1d396[19]),
    .o(al_c81182c));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_79b2ad18 (
    .i(al_55882f9d),
    .o(al_a0e1d396[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a09a83e9 (
    .i(al_a0e1d396[1]),
    .o(al_9b5a4dbd));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5a1feeb5 (
    .i(al_314e2528),
    .o(al_a0e1d396[20]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_631c7f0b (
    .i(al_a0e1d396[20]),
    .o(al_b8da0e9e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_860753e9 (
    .i(al_74f1ae6b),
    .o(al_a0e1d396[21]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_68ddcad7 (
    .i(al_a0e1d396[21]),
    .o(al_fef4ecdb));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_887944ab (
    .i(al_49840bbd),
    .o(al_a0e1d396[22]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c7542061 (
    .i(al_a0e1d396[22]),
    .o(al_796e34c4));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5287ecaf (
    .i(al_fa62f20b),
    .o(al_a0e1d396[23]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1f90a220 (
    .i(al_a0e1d396[23]),
    .o(al_df7aa915));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f8d1aeba (
    .i(al_7da0d957),
    .o(al_a0e1d396[24]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6b9c7c0 (
    .i(al_a0e1d396[24]),
    .o(al_6dc98a03));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_62f6f3e8 (
    .i(al_53b6ba74),
    .o(al_a0e1d396[25]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a241c0bb (
    .i(al_a0e1d396[25]),
    .o(al_80360204));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c3e13c8b (
    .i(al_46888ef2),
    .o(al_a0e1d396[26]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_ca17069 (
    .i(al_a0e1d396[26]),
    .o(al_2bb74c3d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3ca082ca (
    .i(al_8c43abb),
    .o(al_a0e1d396[27]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_696f6a40 (
    .i(al_a0e1d396[27]),
    .o(al_9dcab982));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_e4d44d90 (
    .i(al_89f795c9),
    .o(al_a0e1d396[28]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4bf70c6d (
    .i(al_a0e1d396[28]),
    .o(al_a9490be8));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5ad40da2 (
    .i(al_652cea26),
    .o(al_a0e1d396[29]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_dd711079 (
    .i(al_a0e1d396[29]),
    .o(al_28d8d34d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4fa37ad1 (
    .i(al_267f05f8),
    .o(al_a0e1d396[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_92f37b80 (
    .i(al_a0e1d396[2]),
    .o(al_e6ea44e6));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_17ea5c50 (
    .i(al_2f52bc7e),
    .o(al_a0e1d396[30]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_64e9675c (
    .i(al_a0e1d396[30]),
    .o(al_7cd149c6));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d043dce8 (
    .i(al_14f4e684),
    .o(al_a0e1d396[31]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_bdead46e (
    .i(al_a0e1d396[31]),
    .o(al_b56307ec));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_9db2c7d0 (
    .i(al_1bbf8570),
    .o(al_a0e1d396[32]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_475cb8bb (
    .i(al_a0e1d396[32]),
    .o(al_31be1d74));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ebcacd92 (
    .i(al_59fdd957),
    .o(al_a0e1d396[33]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_96c465eb (
    .i(al_a0e1d396[33]),
    .o(al_cc2e5bcc));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_948e6a74 (
    .i(al_4e23dc54),
    .o(al_a0e1d396[34]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_76086585 (
    .i(al_a0e1d396[34]),
    .o(al_ee615f87));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ca57cba2 (
    .i(al_d79d15f2),
    .o(al_a0e1d396[35]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7bc619f2 (
    .i(al_a0e1d396[35]),
    .o(al_35f768f4));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a00948dd (
    .i(al_e956701b),
    .o(al_a0e1d396[36]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_103d3964 (
    .i(al_a0e1d396[36]),
    .o(al_5e6f3859));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ae509cda (
    .i(al_3ec6ca0b),
    .o(al_a0e1d396[37]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_de1b8068 (
    .i(al_a0e1d396[37]),
    .o(al_2efa36ca));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_fbccc56d (
    .i(al_38793d0),
    .o(al_a0e1d396[38]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e339789a (
    .i(al_a0e1d396[38]),
    .o(al_4708b339));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ec2566a5 (
    .i(al_3ea78ea2),
    .o(al_a0e1d396[39]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7ce09849 (
    .i(al_a0e1d396[39]),
    .o(al_4864d933));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ed69e2d5 (
    .i(al_c600a777),
    .o(al_a0e1d396[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_dc65c0bf (
    .i(al_a0e1d396[3]),
    .o(al_71cac35e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d7981c4a (
    .i(al_c678f752),
    .o(al_a0e1d396[40]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_5765f308 (
    .i(al_a0e1d396[40]),
    .o(al_c3e70575));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_94a774bf (
    .i(al_5f1c8d24),
    .o(al_a0e1d396[41]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_66040bfb (
    .i(al_a0e1d396[41]),
    .o(al_83ebd977));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_84ec6f75 (
    .i(al_ef6225f5),
    .o(al_a0e1d396[42]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2c58ca8 (
    .i(al_a0e1d396[42]),
    .o(al_6bddd01a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a259dffe (
    .i(al_435ecf83),
    .o(al_a0e1d396[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_bb7406c7 (
    .i(al_a0e1d396[4]),
    .o(al_c85cbcb));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1290dc94 (
    .i(al_c802abc3),
    .o(al_a0e1d396[5]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1c976709 (
    .i(al_a0e1d396[5]),
    .o(al_f7c9608b));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_be29f042 (
    .i(al_b6615be3),
    .o(al_a0e1d396[6]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3045e3fa (
    .i(al_a0e1d396[6]),
    .o(al_ac593c94));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b2d944e (
    .i(al_53c183a7),
    .o(al_a0e1d396[7]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_59d31860 (
    .i(al_a0e1d396[7]),
    .o(al_ad58fbc9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ff13d326 (
    .i(al_4b7e1c0f),
    .o(al_a0e1d396[8]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_95f070b2 (
    .i(al_a0e1d396[8]),
    .o(al_3d66f550));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7065aef3 (
    .i(al_228163ab),
    .o(al_a0e1d396[9]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_81b0f088 (
    .i(al_a0e1d396[9]),
    .o(al_12b38499));
  AL_DFF_0 al_cf0fb911 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2d126bfd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5d41495));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a618a9fd (
    .i(al_f5d41495),
    .o(al_d3da8bb7));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7f114e25 (
    .i(al_d3da8bb7),
    .o(al_733c48ff));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_e8e0ed03 (
    .a(al_99c75e01),
    .b(al_5b144427),
    .o(al_2d126bfd[0]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_51e3df6c (
    .a(al_99c75e01),
    .b(al_42d963e6),
    .o(al_2d126bfd[1]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_f17414f3 (
    .a(al_99c75e01),
    .b(al_f1015bac),
    .o(al_2d126bfd[2]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_686f1b42 (
    .a(al_99c75e01),
    .b(al_8cf002a4),
    .o(al_2d126bfd[3]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_de82d5f9 (
    .di(al_19e026e1),
    .raddr(al_620ff4d8[4:0]),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_581e4e41),
    .wclk(al_ef3696df[0]),
    .we(al_733c48ff),
    .rdo(al_b2febcce));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d1fbfce4 (
    .di(al_19e026e1),
    .raddr(al_d23802b0),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_581e4e41),
    .wclk(al_ef3696df[0]),
    .we(al_733c48ff),
    .rdo({open_n270,al_1719553b[0]}));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_4d0875b1 (
    .di(al_3d403a98),
    .raddr(al_8e42692a),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_b16a7f51),
    .wclk(al_ef3696df[0]),
    .we(al_5e87f1a6),
    .rdo({open_n273,al_4caca369[0]}));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3524f5f (
    .di(al_3d403a98),
    .raddr(al_7c49eb0a),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_b16a7f51),
    .wclk(al_ef3696df[0]),
    .we(al_5e87f1a6),
    .rdo({open_n276,al_9681ccaa[0]}));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_a7a834bd (
    .di(al_cc43b80),
    .raddr(al_880139ce),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_f078a0d3),
    .wclk(al_ef3696df[0]),
    .we(al_addcc22),
    .rdo({open_n279,al_b065182c[0]}));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f71b993f (
    .di(al_cc43b80),
    .raddr(al_4d6d3de1),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_f078a0d3),
    .wclk(al_ef3696df[0]),
    .we(al_addcc22),
    .rdo({open_n282,al_1aa44e47[0]}));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ebf43315 (
    .di(al_16418241),
    .raddr(al_8119a127),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_cc30604e),
    .wclk(al_ef3696df[0]),
    .we(al_549369e),
    .rdo({open_n285,al_28515a17[0]}));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_143870ef (
    .di(al_16418241),
    .raddr(al_151512a8),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr(al_cc30604e),
    .wclk(al_ef3696df[0]),
    .we(al_549369e),
    .rdo({open_n288,al_f62892[0]}));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_74a492a9 (
    .i(al_411ed67e),
    .o(al_6b28e3d[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2e06af6b (
    .i(al_6b28e3d[0]),
    .o(al_5e87f1a6));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_e51ebaec (
    .i(al_b00f7d00),
    .o(al_6b28e3d[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_262e690c (
    .i(al_6b28e3d[1]),
    .o(al_addcc22));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_9d200823 (
    .i(al_1342f12a),
    .o(al_6b28e3d[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b934fb5 (
    .i(al_6b28e3d[2]),
    .o(al_549369e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_324314e0 (
    .i(al_4ba727b9),
    .o(al_dfd53060[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_f8d14ee (
    .i(al_dfd53060[0]),
    .o(al_7c49eb0a[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7e58a41e (
    .a(al_511af127[0]),
    .b(al_8e42692a[0]),
    .c(al_42d963e6),
    .o(al_4ba727b9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_90b87609 (
    .i(al_d86483c1),
    .o(al_dfd53060[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_38250343 (
    .i(al_dfd53060[1]),
    .o(al_7c49eb0a[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b4b000a1 (
    .a(al_511af127[1]),
    .b(al_8e42692a[1]),
    .c(al_42d963e6),
    .o(al_d86483c1));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_2d4f43c4 (
    .i(al_5d73fdac),
    .o(al_dfd53060[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b2eb6d2c (
    .i(al_dfd53060[2]),
    .o(al_7c49eb0a[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_10db22a4 (
    .a(al_511af127[2]),
    .b(al_8e42692a[2]),
    .c(al_42d963e6),
    .o(al_5d73fdac));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a56b4d2b (
    .i(al_f4c0ad0d),
    .o(al_dfd53060[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d83a50aa (
    .i(al_dfd53060[3]),
    .o(al_7c49eb0a[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4bc72018 (
    .a(al_511af127[3]),
    .b(al_8e42692a[3]),
    .c(al_42d963e6),
    .o(al_f4c0ad0d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8ab3f0ea (
    .i(al_7b91dfdd),
    .o(al_dfd53060[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_cbb67382 (
    .i(al_dfd53060[4]),
    .o(al_7c49eb0a[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_119e17bb (
    .a(al_511af127[4]),
    .b(al_8e42692a[4]),
    .c(al_42d963e6),
    .o(al_7b91dfdd));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_68b042a8 (
    .i(al_70f2e5bd),
    .o(al_fa928a76[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_143dc9c0 (
    .i(al_fa928a76[0]),
    .o(al_4d6d3de1[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c8eba3f5 (
    .a(al_511af127[0]),
    .b(al_880139ce[0]),
    .c(al_f1015bac),
    .o(al_70f2e5bd));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ce3c060f (
    .i(al_e46ca45e),
    .o(al_fa928a76[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4a9b13d1 (
    .i(al_fa928a76[1]),
    .o(al_4d6d3de1[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_eabeb7b2 (
    .a(al_511af127[1]),
    .b(al_880139ce[1]),
    .c(al_f1015bac),
    .o(al_e46ca45e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_443fe74d (
    .i(al_c77e9fbd),
    .o(al_fa928a76[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7c18cd61 (
    .i(al_fa928a76[2]),
    .o(al_4d6d3de1[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c770b969 (
    .a(al_511af127[2]),
    .b(al_880139ce[2]),
    .c(al_f1015bac),
    .o(al_c77e9fbd));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a6f772b (
    .i(al_62c7fa0b),
    .o(al_fa928a76[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9958d5 (
    .i(al_fa928a76[3]),
    .o(al_4d6d3de1[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a484e346 (
    .a(al_511af127[3]),
    .b(al_880139ce[3]),
    .c(al_f1015bac),
    .o(al_62c7fa0b));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_84051864 (
    .i(al_ff9e30e3),
    .o(al_fa928a76[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3140e10f (
    .i(al_fa928a76[4]),
    .o(al_4d6d3de1[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_bbb47bbe (
    .a(al_511af127[4]),
    .b(al_880139ce[4]),
    .c(al_f1015bac),
    .o(al_ff9e30e3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d13726f (
    .i(al_3cc49650),
    .o(al_7b7033c7[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_134a44af (
    .i(al_7b7033c7[0]),
    .o(al_151512a8[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_138b95b6 (
    .a(al_511af127[0]),
    .b(al_8119a127[0]),
    .c(al_8cf002a4),
    .o(al_3cc49650));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5fb02d1e (
    .i(al_cc952326),
    .o(al_7b7033c7[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b3d38cf8 (
    .i(al_7b7033c7[1]),
    .o(al_151512a8[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1c747aff (
    .a(al_511af127[1]),
    .b(al_8119a127[1]),
    .c(al_8cf002a4),
    .o(al_cc952326));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_fd5ee53d (
    .i(al_2fadb06),
    .o(al_7b7033c7[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b7fab256 (
    .i(al_7b7033c7[2]),
    .o(al_151512a8[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_26033fb (
    .a(al_511af127[2]),
    .b(al_8119a127[2]),
    .c(al_8cf002a4),
    .o(al_2fadb06));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_fe8ce90b (
    .i(al_cf62a4e7),
    .o(al_7b7033c7[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b1944359 (
    .i(al_7b7033c7[3]),
    .o(al_151512a8[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1dd0c7f8 (
    .a(al_511af127[3]),
    .b(al_8119a127[3]),
    .c(al_8cf002a4),
    .o(al_cf62a4e7));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_9976198b (
    .i(al_7fe14516),
    .o(al_7b7033c7[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4d35ef7d (
    .i(al_7b7033c7[4]),
    .o(al_151512a8[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_bd86d352 (
    .a(al_511af127[4]),
    .b(al_8119a127[4]),
    .c(al_8cf002a4),
    .o(al_7fe14516));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5753195a (
    .i(al_a2b915e0),
    .o(al_167833a3[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d236e75d (
    .i(al_167833a3[0]),
    .o(al_b16a7f51[0]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_28ae6a2b (
    .i(al_d0805f59),
    .o(al_167833a3[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_20d8960a (
    .i(al_167833a3[1]),
    .o(al_b16a7f51[1]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ec5adfab (
    .i(al_710215be),
    .o(al_167833a3[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_25ebfc38 (
    .i(al_167833a3[2]),
    .o(al_b16a7f51[2]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8d56a138 (
    .i(al_20e796af),
    .o(al_167833a3[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_60161094 (
    .i(al_167833a3[3]),
    .o(al_b16a7f51[3]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_2526c7d3 (
    .i(al_f567595c),
    .o(al_167833a3[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7655d0a (
    .i(al_167833a3[4]),
    .o(al_b16a7f51[4]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b52402f6 (
    .i(al_d7411c1e),
    .o(al_c85123b0[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_ef92202 (
    .i(al_c85123b0[0]),
    .o(al_f078a0d3[0]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_2a553240 (
    .i(al_4dade993),
    .o(al_c85123b0[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a575a327 (
    .i(al_c85123b0[1]),
    .o(al_f078a0d3[1]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_19e7cf74 (
    .i(al_1ea20fda),
    .o(al_c85123b0[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_5dbc2f9c (
    .i(al_c85123b0[2]),
    .o(al_f078a0d3[2]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8c158e02 (
    .i(al_5f044880),
    .o(al_c85123b0[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3a6086e4 (
    .i(al_c85123b0[3]),
    .o(al_f078a0d3[3]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4d84a202 (
    .i(al_6c6e8c75),
    .o(al_c85123b0[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_574d48c (
    .i(al_c85123b0[4]),
    .o(al_f078a0d3[4]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a58c18db (
    .i(al_b3b929ae),
    .o(al_2b539460[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c3edb597 (
    .i(al_2b539460[0]),
    .o(al_cc30604e[0]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_2327b02c (
    .i(al_cb65ad25),
    .o(al_2b539460[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_f74aeca7 (
    .i(al_2b539460[1]),
    .o(al_cc30604e[1]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c9719b75 (
    .i(al_881adcbc),
    .o(al_2b539460[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d1610486 (
    .i(al_2b539460[2]),
    .o(al_cc30604e[2]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_406c57e8 (
    .i(al_9683b2fb),
    .o(al_2b539460[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_21c8bf34 (
    .i(al_2b539460[3]),
    .o(al_cc30604e[3]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a8c9476 (
    .i(al_7e6b3b5a),
    .o(al_2b539460[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b039196c (
    .i(al_2b539460[4]),
    .o(al_cc30604e[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a25048bd (
    .a(al_511af127[0]),
    .b(al_620ff4d8[0]),
    .c(al_5b144427),
    .o(al_d23802b0[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ff4e6e8e (
    .a(al_511af127[1]),
    .b(al_620ff4d8[1]),
    .c(al_5b144427),
    .o(al_d23802b0[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_abeabe64 (
    .a(al_511af127[2]),
    .b(al_620ff4d8[2]),
    .c(al_5b144427),
    .o(al_d23802b0[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4a23d2f6 (
    .a(al_511af127[3]),
    .b(al_620ff4d8[3]),
    .c(al_5b144427),
    .o(al_d23802b0[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_504a5de5 (
    .a(al_511af127[4]),
    .b(al_620ff4d8[4]),
    .c(al_5b144427),
    .o(al_d23802b0[4]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4df59330 (
    .i(al_2d3877ba),
    .o(al_38d9ed4e[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b40fec65 (
    .i(al_38d9ed4e[0]),
    .o(al_efb91504));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_faf3f745 (
    .a(al_42d963e6),
    .b(al_9681ccaa[0]),
    .o(al_2d3877ba));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_38368104 (
    .i(al_42d963e6),
    .o(al_38d9ed4e[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_65f4fa5 (
    .i(al_38d9ed4e[1]),
    .o(al_60238e88));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_e6f122cc (
    .i(al_691fa5a3),
    .o(al_6c3e2294[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_557e3cb2 (
    .i(al_6c3e2294[0]),
    .o(al_37606c32));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_afb6e3a1 (
    .a(al_f1015bac),
    .b(al_1aa44e47[0]),
    .o(al_691fa5a3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_67232633 (
    .i(al_f1015bac),
    .o(al_6c3e2294[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_8ef7350a (
    .i(al_6c3e2294[1]),
    .o(al_2404250b));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_e70e9912 (
    .i(al_efea142b),
    .o(al_61432edc[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_34e0552e (
    .i(al_61432edc[0]),
    .o(al_5c1ef4c7));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_d81476d (
    .a(al_8cf002a4),
    .b(al_f62892[0]),
    .o(al_efea142b));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7f573647 (
    .i(al_8cf002a4),
    .o(al_61432edc[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3242d24f (
    .i(al_61432edc[1]),
    .o(al_817a8c80));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c4e0a4df (
    .i(al_ac2df9bf),
    .o(al_8f9b22bd[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_8924aa5 (
    .i(al_8f9b22bd[0]),
    .o(al_3d403a98[0]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c965ed82 (
    .i(al_1cb90ce6),
    .o(al_8f9b22bd[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9a2fc03e (
    .i(al_8f9b22bd[1]),
    .o(al_3d403a98[1]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a0a877e7 (
    .i(al_607ca590),
    .o(al_a49512ff[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_328d672d (
    .i(al_a49512ff[0]),
    .o(al_cc43b80[0]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_28f27a39 (
    .i(al_33994c72),
    .o(al_a49512ff[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4b66a177 (
    .i(al_a49512ff[1]),
    .o(al_cc43b80[1]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c9c651fd (
    .i(al_a28bab3a),
    .o(al_d4e10e0d[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d9174046 (
    .i(al_d4e10e0d[0]),
    .o(al_16418241[0]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_54110d5c (
    .i(al_e0914439),
    .o(al_d4e10e0d[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2b3f448f (
    .i(al_d4e10e0d[1]),
    .o(al_16418241[1]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_bb054834 (
    .i(al_48ead91e),
    .o(al_7f5f60b[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b39a805c (
    .i(al_7f5f60b[0]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ba5c95f1 (
    .i(al_a390ad74),
    .o(al_7f5f60b[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_45ab189 (
    .i(al_7f5f60b[1]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_38fa174e (
    .i(al_4c8ccef5),
    .o(al_7f5f60b[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_418eaead (
    .i(al_7f5f60b[2]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_617215b1 (
    .i(al_41c5883),
    .o(al_a51937a3[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_198447b7 (
    .i(al_a51937a3[0]),
    .o(al_2acf9590));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_17546b78 (
    .i(al_361b3557),
    .o(al_a51937a3[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6ed6ccf (
    .i(al_a51937a3[1]),
    .o(al_60b9b0f8));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a28863cb (
    .i(al_54a8a910),
    .o(al_a51937a3[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a34245af (
    .i(al_a51937a3[2]),
    .o(al_f49dc4e0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_26bc7728 (
    .i(al_5f0a94fd),
    .o(al_a51937a3[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_fe042b9e (
    .i(al_a51937a3[3]),
    .o(al_eaa97ed5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_93dd514b (
    .i(al_aa906eb4),
    .o(al_a51937a3[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_12158acb (
    .i(al_a51937a3[4]),
    .o(al_72bfbb1a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_62c423bb (
    .i(al_20745547),
    .o(al_a51937a3[5]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9ca9931a (
    .i(al_a51937a3[5]),
    .o(al_83931c3d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b5a3491 (
    .i(al_8f0f91a1),
    .o(al_a51937a3[6]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_db763812 (
    .i(al_a51937a3[6]),
    .o(al_2117afe8));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c8c7b661 (
    .i(al_7d364519),
    .o(al_a51937a3[7]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_ca8e23aa (
    .i(al_a51937a3[7]),
    .o(al_ebd79caa));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_9db29680 (
    .a(al_162fb89b[0]),
    .b(al_162fb89b[1]),
    .c(al_162fb89b[2]),
    .d(al_162fb89b[3]),
    .e(al_162fb89b[4]),
    .f(al_2acf9590),
    .o(al_50ec922d[0]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_5626e56a (
    .a(al_162fb89b[0]),
    .b(al_162fb89b[1]),
    .c(al_162fb89b[2]),
    .d(al_162fb89b[3]),
    .e(al_162fb89b[4]),
    .f(al_60b9b0f8),
    .o(al_50ec922d[1]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_399da061 (
    .a(al_162fb89b[0]),
    .b(al_162fb89b[1]),
    .c(al_162fb89b[2]),
    .d(al_162fb89b[3]),
    .e(al_162fb89b[4]),
    .f(al_f49dc4e0),
    .o(al_50ec922d[2]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_7f03bcb8 (
    .a(al_162fb89b[0]),
    .b(al_162fb89b[1]),
    .c(al_162fb89b[2]),
    .d(al_162fb89b[3]),
    .e(al_162fb89b[4]),
    .f(al_eaa97ed5),
    .o(al_50ec922d[3]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_eb0be771 (
    .a(al_162fb89b[0]),
    .b(al_162fb89b[1]),
    .c(al_162fb89b[2]),
    .d(al_162fb89b[3]),
    .e(al_162fb89b[4]),
    .f(al_72bfbb1a),
    .o(al_50ec922d[4]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_2cc8f286 (
    .a(al_162fb89b[0]),
    .b(al_162fb89b[1]),
    .c(al_162fb89b[2]),
    .d(al_162fb89b[3]),
    .e(al_162fb89b[4]),
    .f(al_83931c3d),
    .o(al_50ec922d[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_1c9c5fb2 (
    .a(al_162fb89b[0]),
    .b(al_162fb89b[1]),
    .c(al_162fb89b[2]),
    .d(al_162fb89b[3]),
    .e(al_162fb89b[4]),
    .f(al_2117afe8),
    .o(al_50ec922d[6]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*B*A))"),
    .INIT(64'hffffffff80000000))
    al_ca9badd8 (
    .a(al_162fb89b[0]),
    .b(al_162fb89b[1]),
    .c(al_162fb89b[2]),
    .d(al_162fb89b[3]),
    .e(al_162fb89b[4]),
    .f(al_ebd79caa),
    .o(al_50ec922d[7]));
  AL_DFF_0 al_40f2bf99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a90a7b11),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_69b84ba6[2]));
  AL_DFF_0 al_bbf0b61d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2ded3658),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_69b84ba6[3]));
  AL_DFF_0 al_8569b383 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5068e71b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_69b84ba6[4]));
  AL_DFF_0 al_846017e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9ef819de),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_69b84ba6[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_63a48118 (
    .a(ddr_app_rd_data_end),
    .b(al_70117344),
    .o(al_6b872c5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hdffffffffffffffb))
    al_b9989ab1 (
    .a(al_a7c937ec),
    .b(al_6b872c5),
    .c(al_69b84ba6[0]),
    .d(al_69b84ba6[1]),
    .e(al_69b84ba6[2]),
    .f(al_69b84ba6[3]),
    .o(al_58e4bd8e));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_526c6e38 (
    .a(al_69b84ba6[0]),
    .b(al_69b84ba6[1]),
    .c(al_69b84ba6[2]),
    .d(al_69b84ba6[3]),
    .e(al_69b84ba6[4]),
    .o(al_fdaccc20));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_4841938b (
    .a(al_58e4bd8e),
    .b(al_6db5b9d2),
    .c(al_69b84ba6[4]),
    .o(al_5068e71b));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D@B@A))"),
    .INIT(16'h0906))
    al_65baab27 (
    .a(al_a7c937ec),
    .b(al_6b872c5),
    .c(al_6db5b9d2),
    .d(al_69b84ba6[0]),
    .o(al_5ace851));
  AL_MAP_LUT6 #(
    .EQN("(~C*(F@(~(A)*B*~(D)*~(E)+A*~(B)*D*E)))"),
    .INIT(64'h0d0f0f0b02000004))
    al_7143e38a (
    .a(al_a7c937ec),
    .b(al_6b872c5),
    .c(al_6db5b9d2),
    .d(al_69b84ba6[0]),
    .e(al_69b84ba6[1]),
    .f(al_69b84ba6[2]),
    .o(al_a90a7b11));
  AL_MAP_LUT6 #(
    .EQN("(F@(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h20000004dffffffb))
    al_ed9f39e2 (
    .a(al_a7c937ec),
    .b(al_6b872c5),
    .c(al_69b84ba6[0]),
    .d(al_69b84ba6[1]),
    .e(al_69b84ba6[2]),
    .f(al_69b84ba6[3]),
    .o(al_ce84f7a6));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_7b647426 (
    .a(al_ce84f7a6),
    .b(al_6db5b9d2),
    .o(al_2ded3658));
  AL_MAP_LUT5 #(
    .EQN("(~C*(E@(~(A)*B*~(D)+A*~(B)*D)))"),
    .INIT(32'h0d0b0204))
    al_40fa031e (
    .a(al_a7c937ec),
    .b(al_6b872c5),
    .c(al_6db5b9d2),
    .d(al_69b84ba6[0]),
    .e(al_69b84ba6[1]),
    .o(al_e825eb09));
  AL_MAP_LUT6 #(
    .EQN("(~E*(F@(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*B*C*D)))"),
    .INIT(64'h0000bb5f000044a0))
    al_9e24ae0 (
    .a(al_a7c937ec),
    .b(al_fdaccc20),
    .c(al_71fc1ad7),
    .d(al_6b872c5),
    .e(al_6db5b9d2),
    .f(al_69b84ba6[5]),
    .o(al_9ef819de));
  AL_DFF_0 al_afbaa783 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5ace851),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_69b84ba6[0]));
  AL_DFF_0 al_4b7f4083 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e825eb09),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_69b84ba6[1]));
  AL_DFF_0 al_3d79ca89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9d23d003),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_100c2219[2]));
  AL_DFF_0 al_f57d003 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a12892b0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_100c2219[3]));
  AL_DFF_0 al_ef4af5b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ddd2e3de),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_100c2219[4]));
  AL_DFF_0 al_199c458b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_de2b5681),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_100c2219[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_98e0e4a5 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_100c2219[0]),
    .e(al_100c2219[1]),
    .f(al_100c2219[2]),
    .o(al_fd874a49));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_263b0aca (
    .a(al_fd874a49),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_100c2219[3]),
    .f(al_100c2219[4]),
    .o(al_3728ce00));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_7b9bde12 (
    .a(al_3728ce00),
    .b(al_100c2219[5]),
    .c(al_df90085e),
    .d(al_4caca369[0]),
    .o(al_4830d0fa));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_c3fdcd73 (
    .a(al_4830d0fa),
    .b(al_100c2219[0]),
    .c(al_100c2219[1]),
    .o(al_b0eff5ca));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_4b39897b (
    .a(al_b0eff5ca),
    .b(al_6db5b9d2),
    .c(al_100c2219[2]),
    .d(al_100c2219[3]),
    .e(al_100c2219[4]),
    .o(al_ddd2e3de));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_409c6074 (
    .a(al_b0eff5ca),
    .b(al_6db5b9d2),
    .c(al_100c2219[2]),
    .d(al_100c2219[3]),
    .o(al_a12892b0));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_32d7dd2 (
    .a(al_4830d0fa),
    .b(al_6db5b9d2),
    .c(al_100c2219[0]),
    .o(al_11041b8b));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_655dad73 (
    .a(al_4830d0fa),
    .b(al_6db5b9d2),
    .c(al_100c2219[0]),
    .d(al_100c2219[1]),
    .o(al_fe081845));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_d15d839 (
    .a(al_b0eff5ca),
    .b(al_6db5b9d2),
    .c(al_100c2219[2]),
    .o(al_9d23d003));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_9789db1 (
    .a(al_b0eff5ca),
    .b(al_6db5b9d2),
    .c(al_100c2219[2]),
    .d(al_100c2219[3]),
    .e(al_100c2219[4]),
    .f(al_100c2219[5]),
    .o(al_de2b5681));
  AL_DFF_0 al_20ecad94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_11041b8b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_100c2219[0]));
  AL_DFF_0 al_d55b202d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fe081845),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_100c2219[1]));
  AL_DFF_0 al_4a741210 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c6d66579),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2d22d77a[2]));
  AL_DFF_0 al_825dd1b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a9ffc103),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2d22d77a[3]));
  AL_DFF_0 al_ea187dfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7ee48c14),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2d22d77a[4]));
  AL_DFF_0 al_59d9f46b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2599c30),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2d22d77a[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_239852e6 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_2d22d77a[0]),
    .e(al_2d22d77a[1]),
    .f(al_2d22d77a[2]),
    .o(al_5679c3a4));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_ecf1dc58 (
    .a(al_5679c3a4),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_2d22d77a[3]),
    .f(al_2d22d77a[4]),
    .o(al_a6167193));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_15189b3a (
    .a(al_a6167193),
    .b(al_2d22d77a[5]),
    .c(al_72ab91cb),
    .d(al_b065182c[0]),
    .o(al_1b9ef62a));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_58110640 (
    .a(al_1b9ef62a),
    .b(al_2d22d77a[0]),
    .c(al_2d22d77a[1]),
    .o(al_9ab94adf));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_cdd913 (
    .a(al_9ab94adf),
    .b(al_6db5b9d2),
    .c(al_2d22d77a[2]),
    .d(al_2d22d77a[3]),
    .e(al_2d22d77a[4]),
    .o(al_7ee48c14));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_c5e951db (
    .a(al_9ab94adf),
    .b(al_6db5b9d2),
    .c(al_2d22d77a[2]),
    .d(al_2d22d77a[3]),
    .o(al_a9ffc103));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_fa696e25 (
    .a(al_1b9ef62a),
    .b(al_6db5b9d2),
    .c(al_2d22d77a[0]),
    .o(al_fd64f6c3));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_55443cc4 (
    .a(al_1b9ef62a),
    .b(al_6db5b9d2),
    .c(al_2d22d77a[0]),
    .d(al_2d22d77a[1]),
    .o(al_d3947eeb));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_1767ba8a (
    .a(al_9ab94adf),
    .b(al_6db5b9d2),
    .c(al_2d22d77a[2]),
    .o(al_c6d66579));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_52b9ba8b (
    .a(al_9ab94adf),
    .b(al_6db5b9d2),
    .c(al_2d22d77a[2]),
    .d(al_2d22d77a[3]),
    .e(al_2d22d77a[4]),
    .f(al_2d22d77a[5]),
    .o(al_2599c30));
  AL_DFF_0 al_cb6646a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd64f6c3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2d22d77a[0]));
  AL_DFF_0 al_3b8b40b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d3947eeb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2d22d77a[1]));
  AL_DFF_0 al_e4607c54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dd2698f4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8af537d6[2]));
  AL_DFF_0 al_9f02e80c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_793e445),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8af537d6[3]));
  AL_DFF_0 al_e99a0f98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_858348d9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8af537d6[4]));
  AL_DFF_0 al_bf3fe9b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e2481062),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8af537d6[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_a5c08336 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_8af537d6[0]),
    .e(al_8af537d6[1]),
    .f(al_8af537d6[2]),
    .o(al_ba7f7c4));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_4b1c8314 (
    .a(al_ba7f7c4),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_8af537d6[3]),
    .f(al_8af537d6[4]),
    .o(al_3310bf9b));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_6e176690 (
    .a(al_3310bf9b),
    .b(al_8af537d6[5]),
    .c(al_c9d182cf),
    .d(al_28515a17[0]),
    .o(al_3f0f44a5));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_1fa6426e (
    .a(al_3f0f44a5),
    .b(al_8af537d6[0]),
    .c(al_8af537d6[1]),
    .o(al_ee9d432a));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_18a713 (
    .a(al_ee9d432a),
    .b(al_6db5b9d2),
    .c(al_8af537d6[2]),
    .d(al_8af537d6[3]),
    .e(al_8af537d6[4]),
    .o(al_858348d9));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_3157d45f (
    .a(al_ee9d432a),
    .b(al_6db5b9d2),
    .c(al_8af537d6[2]),
    .d(al_8af537d6[3]),
    .o(al_793e445));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_bc56a49a (
    .a(al_3f0f44a5),
    .b(al_6db5b9d2),
    .c(al_8af537d6[0]),
    .o(al_799ff6e6));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_8fedbd10 (
    .a(al_3f0f44a5),
    .b(al_6db5b9d2),
    .c(al_8af537d6[0]),
    .d(al_8af537d6[1]),
    .o(al_eb0a7105));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_44ea104c (
    .a(al_ee9d432a),
    .b(al_6db5b9d2),
    .c(al_8af537d6[2]),
    .o(al_dd2698f4));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_51551176 (
    .a(al_ee9d432a),
    .b(al_6db5b9d2),
    .c(al_8af537d6[2]),
    .d(al_8af537d6[3]),
    .e(al_8af537d6[4]),
    .f(al_8af537d6[5]),
    .o(al_e2481062));
  AL_DFF_0 al_dbadc377 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_799ff6e6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8af537d6[0]));
  AL_DFF_0 al_dffec844 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eb0a7105),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8af537d6[1]));
  AL_DFF_0 al_e0ac02b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ce170fdf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_175608a7[2]));
  AL_DFF_0 al_2259d010 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_19a0944b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_175608a7[3]));
  AL_DFF_0 al_cd316823 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eaa78f2d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_175608a7[4]));
  AL_DFF_0 al_3147a603 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b7614e0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_175608a7[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_ee3d7230 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_175608a7[0]),
    .e(al_175608a7[1]),
    .f(al_175608a7[2]),
    .o(al_79846c19));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_486b320a (
    .a(al_79846c19),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_175608a7[3]),
    .f(al_175608a7[4]),
    .o(al_af74714f));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_66e51679 (
    .a(al_af74714f),
    .b(al_175608a7[5]),
    .c(al_4f9aa153),
    .d(al_4caca369[0]),
    .o(al_ab431a20));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_7adc2716 (
    .a(al_ab431a20),
    .b(al_175608a7[0]),
    .c(al_175608a7[1]),
    .o(al_f2d75fa6));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_9eca9a32 (
    .a(al_f2d75fa6),
    .b(al_6db5b9d2),
    .c(al_175608a7[2]),
    .d(al_175608a7[3]),
    .e(al_175608a7[4]),
    .o(al_eaa78f2d));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_269ac1ac (
    .a(al_f2d75fa6),
    .b(al_6db5b9d2),
    .c(al_175608a7[2]),
    .d(al_175608a7[3]),
    .o(al_19a0944b));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_b5c5cffb (
    .a(al_ab431a20),
    .b(al_6db5b9d2),
    .c(al_175608a7[0]),
    .o(al_2eed0a97));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_5195e48a (
    .a(al_ab431a20),
    .b(al_6db5b9d2),
    .c(al_175608a7[0]),
    .d(al_175608a7[1]),
    .o(al_264acb9b));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_e8c5c460 (
    .a(al_f2d75fa6),
    .b(al_6db5b9d2),
    .c(al_175608a7[2]),
    .o(al_ce170fdf));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_68dfdcd4 (
    .a(al_f2d75fa6),
    .b(al_6db5b9d2),
    .c(al_175608a7[2]),
    .d(al_175608a7[3]),
    .e(al_175608a7[4]),
    .f(al_175608a7[5]),
    .o(al_7b7614e0));
  AL_DFF_0 al_cbddfbe6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2eed0a97),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_175608a7[0]));
  AL_DFF_0 al_22869c9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_264acb9b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_175608a7[1]));
  AL_DFF_0 al_de5cb1e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a735e2bc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5e6b3f5[2]));
  AL_DFF_0 al_5f8bae77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_99214f52),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5e6b3f5[3]));
  AL_DFF_0 al_ed51aaa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b58c5a7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5e6b3f5[4]));
  AL_DFF_0 al_4086ba01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b578c72c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5e6b3f5[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_7155390d (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_f5e6b3f5[0]),
    .e(al_f5e6b3f5[1]),
    .f(al_f5e6b3f5[2]),
    .o(al_42d1f999));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_47a9478f (
    .a(al_42d1f999),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_f5e6b3f5[3]),
    .f(al_f5e6b3f5[4]),
    .o(al_8091f068));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_87ccee22 (
    .a(al_8091f068),
    .b(al_f5e6b3f5[5]),
    .c(al_d4c409ba),
    .d(al_b065182c[0]),
    .o(al_f0eae58e));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_282e0141 (
    .a(al_f0eae58e),
    .b(al_f5e6b3f5[0]),
    .c(al_f5e6b3f5[1]),
    .d(al_f5e6b3f5[2]),
    .e(al_f5e6b3f5[3]),
    .f(al_f5e6b3f5[4]),
    .o(al_ed6ca683));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_eaf52dbb (
    .a(al_f0eae58e),
    .b(al_f5e6b3f5[0]),
    .c(al_f5e6b3f5[1]),
    .d(al_f5e6b3f5[2]),
    .e(al_f5e6b3f5[3]),
    .f(al_f5e6b3f5[4]),
    .o(al_ab2d2d18));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_1d8f9424 (
    .a(al_ab2d2d18),
    .b(al_6db5b9d2),
    .o(al_5b58c5a7));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_4a67c964 (
    .a(al_f0eae58e),
    .b(al_6db5b9d2),
    .c(al_f5e6b3f5[0]),
    .d(al_f5e6b3f5[1]),
    .e(al_f5e6b3f5[2]),
    .f(al_f5e6b3f5[3]),
    .o(al_99214f52));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_29d17576 (
    .a(al_f0eae58e),
    .b(al_6db5b9d2),
    .c(al_f5e6b3f5[0]),
    .o(al_beea7df8));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_a0cccac8 (
    .a(al_f0eae58e),
    .b(al_6db5b9d2),
    .c(al_f5e6b3f5[0]),
    .d(al_f5e6b3f5[1]),
    .o(al_6694e9cf));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_5c7d158c (
    .a(al_f0eae58e),
    .b(al_6db5b9d2),
    .c(al_f5e6b3f5[0]),
    .d(al_f5e6b3f5[1]),
    .e(al_f5e6b3f5[2]),
    .o(al_a735e2bc));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_ea28cd73 (
    .a(al_ed6ca683),
    .b(al_6db5b9d2),
    .c(al_f5e6b3f5[5]),
    .o(al_b578c72c));
  AL_DFF_0 al_dc184b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_beea7df8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5e6b3f5[0]));
  AL_DFF_0 al_6cc08305 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6694e9cf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5e6b3f5[1]));
  AL_DFF_0 al_bf1fb1a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7ee9bd9c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_abd25e4c[2]));
  AL_DFF_0 al_25d73bf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b5e551b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_abd25e4c[3]));
  AL_DFF_0 al_77e33905 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3613b64a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_abd25e4c[4]));
  AL_DFF_0 al_e99ae9c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1c42289),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_abd25e4c[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_92732f31 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_abd25e4c[0]),
    .e(al_abd25e4c[1]),
    .f(al_abd25e4c[2]),
    .o(al_2b594476));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_e6052fa0 (
    .a(al_2b594476),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_abd25e4c[3]),
    .f(al_abd25e4c[4]),
    .o(al_3bfb38e8));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_fffeb417 (
    .a(al_3bfb38e8),
    .b(al_abd25e4c[5]),
    .c(al_e2476620),
    .d(al_b065182c[0]),
    .o(al_41ff936b));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_955c4a9c (
    .a(al_41ff936b),
    .b(al_abd25e4c[0]),
    .c(al_abd25e4c[1]),
    .o(al_97559555));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_b36f1168 (
    .a(al_97559555),
    .b(al_6db5b9d2),
    .c(al_abd25e4c[2]),
    .d(al_abd25e4c[3]),
    .e(al_abd25e4c[4]),
    .o(al_3613b64a));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_b90a3e78 (
    .a(al_97559555),
    .b(al_6db5b9d2),
    .c(al_abd25e4c[2]),
    .d(al_abd25e4c[3]),
    .o(al_7b5e551b));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_271baad2 (
    .a(al_41ff936b),
    .b(al_6db5b9d2),
    .c(al_abd25e4c[0]),
    .o(al_366699aa));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_3245a89 (
    .a(al_41ff936b),
    .b(al_6db5b9d2),
    .c(al_abd25e4c[0]),
    .d(al_abd25e4c[1]),
    .o(al_cffc4db7));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_e8bc7094 (
    .a(al_97559555),
    .b(al_6db5b9d2),
    .c(al_abd25e4c[2]),
    .o(al_7ee9bd9c));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_11a333e5 (
    .a(al_97559555),
    .b(al_6db5b9d2),
    .c(al_abd25e4c[2]),
    .d(al_abd25e4c[3]),
    .e(al_abd25e4c[4]),
    .f(al_abd25e4c[5]),
    .o(al_1c42289));
  AL_DFF_0 al_29f0dd2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_366699aa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_abd25e4c[0]));
  AL_DFF_0 al_30a6c88e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cffc4db7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_abd25e4c[1]));
  AL_DFF_0 al_9c560cd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_754cb61b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9cdd3a01[2]));
  AL_DFF_0 al_31bd81bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8f668693),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9cdd3a01[3]));
  AL_DFF_0 al_79f019db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_815d1ad6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9cdd3a01[4]));
  AL_DFF_0 al_6cf7cdb6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_757240b3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9cdd3a01[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_5402eb78 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_9cdd3a01[0]),
    .e(al_9cdd3a01[1]),
    .f(al_9cdd3a01[2]),
    .o(al_1dbc8101));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_3ecc1925 (
    .a(al_1dbc8101),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_9cdd3a01[3]),
    .f(al_9cdd3a01[4]),
    .o(al_ad24301));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_2263bb64 (
    .a(al_ad24301),
    .b(al_9cdd3a01[5]),
    .c(al_24944e5c),
    .d(al_28515a17[0]),
    .o(al_2d8e01f3));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_ded62199 (
    .a(al_2d8e01f3),
    .b(al_9cdd3a01[0]),
    .c(al_9cdd3a01[1]),
    .o(al_8825809e));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_f581108f (
    .a(al_8825809e),
    .b(al_6db5b9d2),
    .c(al_9cdd3a01[2]),
    .d(al_9cdd3a01[3]),
    .e(al_9cdd3a01[4]),
    .o(al_815d1ad6));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_7cd1ceb6 (
    .a(al_8825809e),
    .b(al_6db5b9d2),
    .c(al_9cdd3a01[2]),
    .d(al_9cdd3a01[3]),
    .o(al_8f668693));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_b36e4eaf (
    .a(al_2d8e01f3),
    .b(al_6db5b9d2),
    .c(al_9cdd3a01[0]),
    .o(al_613310ab));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_3f01565 (
    .a(al_2d8e01f3),
    .b(al_6db5b9d2),
    .c(al_9cdd3a01[0]),
    .d(al_9cdd3a01[1]),
    .o(al_821df217));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_befe395e (
    .a(al_8825809e),
    .b(al_6db5b9d2),
    .c(al_9cdd3a01[2]),
    .o(al_754cb61b));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_337e4a35 (
    .a(al_8825809e),
    .b(al_6db5b9d2),
    .c(al_9cdd3a01[2]),
    .d(al_9cdd3a01[3]),
    .e(al_9cdd3a01[4]),
    .f(al_9cdd3a01[5]),
    .o(al_757240b3));
  AL_DFF_0 al_9244397c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_613310ab),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9cdd3a01[0]));
  AL_DFF_0 al_599010ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_821df217),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9cdd3a01[1]));
  AL_DFF_0 al_2fa9d235 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ce8339bf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ef04c8[2]));
  AL_DFF_0 al_3975ed4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_18a07add),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ef04c8[3]));
  AL_DFF_0 al_e6aec060 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3339143),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ef04c8[4]));
  AL_DFF_0 al_5a668e8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e7e914bb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ef04c8[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_a5c478bd (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_55ef04c8[0]),
    .e(al_55ef04c8[1]),
    .f(al_55ef04c8[2]),
    .o(al_1506e6b3));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_e1c97aa (
    .a(al_1506e6b3),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_55ef04c8[3]),
    .f(al_55ef04c8[4]),
    .o(al_a4c76fab));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_2596c8cd (
    .a(al_a4c76fab),
    .b(al_55ef04c8[5]),
    .c(al_e2f3bed2),
    .d(al_4caca369[0]),
    .o(al_32c129b3));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_595c6788 (
    .a(al_32c129b3),
    .b(al_55ef04c8[0]),
    .c(al_55ef04c8[1]),
    .o(al_f5ca45d2));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_59284373 (
    .a(al_f5ca45d2),
    .b(al_6db5b9d2),
    .c(al_55ef04c8[2]),
    .d(al_55ef04c8[3]),
    .e(al_55ef04c8[4]),
    .o(al_c3339143));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_4a0723e3 (
    .a(al_f5ca45d2),
    .b(al_6db5b9d2),
    .c(al_55ef04c8[2]),
    .d(al_55ef04c8[3]),
    .o(al_18a07add));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_11a79e65 (
    .a(al_32c129b3),
    .b(al_6db5b9d2),
    .c(al_55ef04c8[0]),
    .o(al_90caa0c7));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_5868a0c3 (
    .a(al_32c129b3),
    .b(al_6db5b9d2),
    .c(al_55ef04c8[0]),
    .d(al_55ef04c8[1]),
    .o(al_1dd9faa9));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_6808521e (
    .a(al_f5ca45d2),
    .b(al_6db5b9d2),
    .c(al_55ef04c8[2]),
    .o(al_ce8339bf));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_6cc34edc (
    .a(al_f5ca45d2),
    .b(al_6db5b9d2),
    .c(al_55ef04c8[2]),
    .d(al_55ef04c8[3]),
    .e(al_55ef04c8[4]),
    .f(al_55ef04c8[5]),
    .o(al_e7e914bb));
  AL_DFF_0 al_3e984f64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_90caa0c7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ef04c8[0]));
  AL_DFF_0 al_aecf70d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1dd9faa9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55ef04c8[1]));
  AL_DFF_0 al_5a0aa375 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4053f9a0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_384dd51d[2]));
  AL_DFF_0 al_4aea4538 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_36161b0f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_384dd51d[3]));
  AL_DFF_0 al_2a788094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2775bd20),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_384dd51d[4]));
  AL_DFF_0 al_cbd8f476 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_290f1dfa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_384dd51d[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_5c11cc84 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_384dd51d[0]),
    .e(al_384dd51d[1]),
    .f(al_384dd51d[2]),
    .o(al_65787e3f));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_a0e7fbb1 (
    .a(al_65787e3f),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_384dd51d[3]),
    .f(al_384dd51d[4]),
    .o(al_f07cc0e));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_2d9787aa (
    .a(al_f07cc0e),
    .b(al_384dd51d[5]),
    .c(al_6db10ea9),
    .d(al_b065182c[0]),
    .o(al_57d1b933));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_2949a527 (
    .a(al_57d1b933),
    .b(al_384dd51d[0]),
    .c(al_384dd51d[1]),
    .o(al_45e32f1a));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_5700a076 (
    .a(al_45e32f1a),
    .b(al_6db5b9d2),
    .c(al_384dd51d[2]),
    .d(al_384dd51d[3]),
    .e(al_384dd51d[4]),
    .o(al_2775bd20));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_795aea18 (
    .a(al_45e32f1a),
    .b(al_6db5b9d2),
    .c(al_384dd51d[2]),
    .d(al_384dd51d[3]),
    .o(al_36161b0f));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_49ae4b23 (
    .a(al_57d1b933),
    .b(al_6db5b9d2),
    .c(al_384dd51d[0]),
    .o(al_60141953));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_d139227 (
    .a(al_57d1b933),
    .b(al_6db5b9d2),
    .c(al_384dd51d[0]),
    .d(al_384dd51d[1]),
    .o(al_cf94ebc3));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_aec3211f (
    .a(al_45e32f1a),
    .b(al_6db5b9d2),
    .c(al_384dd51d[2]),
    .o(al_4053f9a0));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_9d2b775e (
    .a(al_45e32f1a),
    .b(al_6db5b9d2),
    .c(al_384dd51d[2]),
    .d(al_384dd51d[3]),
    .e(al_384dd51d[4]),
    .f(al_384dd51d[5]),
    .o(al_290f1dfa));
  AL_DFF_0 al_8befa6dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_60141953),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_384dd51d[0]));
  AL_DFF_0 al_93370ce0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf94ebc3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_384dd51d[1]));
  AL_DFF_0 al_11744c4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6f3de2dc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_269b6545[2]));
  AL_DFF_0 al_de6add1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_60fd4192),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_269b6545[3]));
  AL_DFF_0 al_d46cf424 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f2987856),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_269b6545[4]));
  AL_DFF_0 al_2f741c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba1ded0d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_269b6545[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_e514c62c (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_269b6545[0]),
    .e(al_269b6545[1]),
    .f(al_269b6545[2]),
    .o(al_4b87de86));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_8fc0eb4b (
    .a(al_4b87de86),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_269b6545[3]),
    .f(al_269b6545[4]),
    .o(al_d8d52ddc));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_3d39ea02 (
    .a(al_d8d52ddc),
    .b(al_269b6545[5]),
    .c(al_7bbb36d3),
    .d(al_28515a17[0]),
    .o(al_32460991));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_afc2f8e9 (
    .a(al_32460991),
    .b(al_269b6545[0]),
    .c(al_269b6545[1]),
    .o(al_a92f34f8));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_82978121 (
    .a(al_a92f34f8),
    .b(al_6db5b9d2),
    .c(al_269b6545[2]),
    .d(al_269b6545[3]),
    .e(al_269b6545[4]),
    .o(al_f2987856));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_26a05696 (
    .a(al_a92f34f8),
    .b(al_6db5b9d2),
    .c(al_269b6545[2]),
    .d(al_269b6545[3]),
    .o(al_60fd4192));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_8312af6a (
    .a(al_32460991),
    .b(al_6db5b9d2),
    .c(al_269b6545[0]),
    .o(al_f3161340));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_7e3655e4 (
    .a(al_32460991),
    .b(al_6db5b9d2),
    .c(al_269b6545[0]),
    .d(al_269b6545[1]),
    .o(al_2570708b));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_bbe34a94 (
    .a(al_a92f34f8),
    .b(al_6db5b9d2),
    .c(al_269b6545[2]),
    .o(al_6f3de2dc));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_c9479bfe (
    .a(al_a92f34f8),
    .b(al_6db5b9d2),
    .c(al_269b6545[2]),
    .d(al_269b6545[3]),
    .e(al_269b6545[4]),
    .f(al_269b6545[5]),
    .o(al_ba1ded0d));
  AL_DFF_0 al_fcbc1f29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3161340),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_269b6545[0]));
  AL_DFF_0 al_687fbcb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2570708b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_269b6545[1]));
  AL_DFF_0 al_6a30f22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c1ffe8c),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_4e8fb619));
  AL_DFF_0 al_42ad49c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2db7ae9f),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_fd6a3ba4));
  AL_DFF_0 al_cd04395f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_adc73f46),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_b3cfcb5e));
  AL_DFF_0 al_f3ec7457 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_99dca23),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_9a7b3b80));
  AL_DFF_0 al_1a81d355 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c9258181),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_430dd919[2]));
  AL_DFF_0 al_20ede004 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_478aa8b9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_430dd919[3]));
  AL_DFF_0 al_fd688ee1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_94a7a40),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_430dd919[4]));
  AL_DFF_0 al_d23f01ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2a63dd17),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_430dd919[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_45148187 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_430dd919[0]),
    .e(al_430dd919[1]),
    .f(al_430dd919[2]),
    .o(al_1081a2ca));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_a43fc5de (
    .a(al_1081a2ca),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_430dd919[3]),
    .f(al_430dd919[4]),
    .o(al_b49bcb3));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_59b03cfa (
    .a(al_b49bcb3),
    .b(al_430dd919[5]),
    .c(al_8d8df5a3),
    .d(al_4caca369[0]),
    .o(al_4704250e));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_740cce06 (
    .a(al_4704250e),
    .b(al_430dd919[0]),
    .c(al_430dd919[1]),
    .d(al_430dd919[2]),
    .e(al_430dd919[3]),
    .f(al_430dd919[4]),
    .o(al_432975cc));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_6d415a55 (
    .a(al_4704250e),
    .b(al_430dd919[0]),
    .c(al_430dd919[1]),
    .d(al_430dd919[2]),
    .e(al_430dd919[3]),
    .f(al_430dd919[4]),
    .o(al_6c74032f));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_bbdf34f0 (
    .a(al_6c74032f),
    .b(al_6db5b9d2),
    .o(al_94a7a40));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_4f3980e (
    .a(al_4704250e),
    .b(al_6db5b9d2),
    .c(al_430dd919[0]),
    .d(al_430dd919[1]),
    .e(al_430dd919[2]),
    .f(al_430dd919[3]),
    .o(al_478aa8b9));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_4fece155 (
    .a(al_4704250e),
    .b(al_6db5b9d2),
    .c(al_430dd919[0]),
    .o(al_a91a268));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_d5d64d92 (
    .a(al_4704250e),
    .b(al_6db5b9d2),
    .c(al_430dd919[0]),
    .d(al_430dd919[1]),
    .o(al_14184769));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_3e584f21 (
    .a(al_4704250e),
    .b(al_6db5b9d2),
    .c(al_430dd919[0]),
    .d(al_430dd919[1]),
    .e(al_430dd919[2]),
    .o(al_c9258181));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_450afab7 (
    .a(al_432975cc),
    .b(al_6db5b9d2),
    .c(al_430dd919[5]),
    .o(al_2a63dd17));
  AL_DFF_0 al_695fb698 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a91a268),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_430dd919[0]));
  AL_DFF_0 al_de389769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_14184769),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_430dd919[1]));
  AL_DFF_0 al_c6d6691d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dc492d87),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c6ba19f[2]));
  AL_DFF_0 al_1d8628bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c37042bd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c6ba19f[3]));
  AL_DFF_0 al_bcc1ad9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_944bd830),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c6ba19f[4]));
  AL_DFF_0 al_bc2f7680 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3624cfe0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c6ba19f[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_9868473f (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_5c6ba19f[0]),
    .e(al_5c6ba19f[1]),
    .f(al_5c6ba19f[2]),
    .o(al_3d1dbb20));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_b7d9a750 (
    .a(al_3d1dbb20),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_5c6ba19f[3]),
    .f(al_5c6ba19f[4]),
    .o(al_312b2dca));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_ded9465b (
    .a(al_312b2dca),
    .b(al_5c6ba19f[5]),
    .c(al_2fc8b96e),
    .d(al_b065182c[0]),
    .o(al_12dd86af));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_3c677ae9 (
    .a(al_12dd86af),
    .b(al_5c6ba19f[0]),
    .c(al_5c6ba19f[1]),
    .o(al_189dc8c0));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_4c4de5c7 (
    .a(al_189dc8c0),
    .b(al_6db5b9d2),
    .c(al_5c6ba19f[2]),
    .d(al_5c6ba19f[3]),
    .e(al_5c6ba19f[4]),
    .o(al_944bd830));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_352be84e (
    .a(al_189dc8c0),
    .b(al_6db5b9d2),
    .c(al_5c6ba19f[2]),
    .d(al_5c6ba19f[3]),
    .o(al_c37042bd));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_9ef59b90 (
    .a(al_12dd86af),
    .b(al_6db5b9d2),
    .c(al_5c6ba19f[0]),
    .o(al_dfa5ff6c));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_8fd52bb0 (
    .a(al_12dd86af),
    .b(al_6db5b9d2),
    .c(al_5c6ba19f[0]),
    .d(al_5c6ba19f[1]),
    .o(al_d211a035));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_fdf4139b (
    .a(al_189dc8c0),
    .b(al_6db5b9d2),
    .c(al_5c6ba19f[2]),
    .o(al_dc492d87));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_80690372 (
    .a(al_189dc8c0),
    .b(al_6db5b9d2),
    .c(al_5c6ba19f[2]),
    .d(al_5c6ba19f[3]),
    .e(al_5c6ba19f[4]),
    .f(al_5c6ba19f[5]),
    .o(al_3624cfe0));
  AL_DFF_0 al_d867aa3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dfa5ff6c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c6ba19f[0]));
  AL_DFF_0 al_e5d5d654 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d211a035),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c6ba19f[1]));
  AL_DFF_0 al_42c1b4dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_34c94edb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f6bae56[2]));
  AL_DFF_0 al_ce29f787 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4ca26c83),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f6bae56[3]));
  AL_DFF_0 al_5721cbc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1a3a4ed7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f6bae56[4]));
  AL_DFF_0 al_98bd5317 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f60ec0d5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f6bae56[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_6253f13c (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_4f6bae56[0]),
    .e(al_4f6bae56[1]),
    .f(al_4f6bae56[2]),
    .o(al_b2e217b));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_b5a57520 (
    .a(al_b2e217b),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_4f6bae56[3]),
    .f(al_4f6bae56[4]),
    .o(al_9b71a4e4));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_3ceb6bda (
    .a(al_9b71a4e4),
    .b(al_4f6bae56[5]),
    .c(al_d27a1279),
    .d(al_28515a17[0]),
    .o(al_df5418e9));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_5b210670 (
    .a(al_df5418e9),
    .b(al_4f6bae56[0]),
    .c(al_4f6bae56[1]),
    .o(al_83ae9a40));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_a8b3a6b4 (
    .a(al_83ae9a40),
    .b(al_6db5b9d2),
    .c(al_4f6bae56[2]),
    .d(al_4f6bae56[3]),
    .e(al_4f6bae56[4]),
    .o(al_1a3a4ed7));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_e4a2a513 (
    .a(al_83ae9a40),
    .b(al_6db5b9d2),
    .c(al_4f6bae56[2]),
    .d(al_4f6bae56[3]),
    .o(al_4ca26c83));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_321b3ea6 (
    .a(al_df5418e9),
    .b(al_6db5b9d2),
    .c(al_4f6bae56[0]),
    .o(al_9609a6f5));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_58eb89c4 (
    .a(al_df5418e9),
    .b(al_6db5b9d2),
    .c(al_4f6bae56[0]),
    .d(al_4f6bae56[1]),
    .o(al_bf0c650));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_d231968d (
    .a(al_83ae9a40),
    .b(al_6db5b9d2),
    .c(al_4f6bae56[2]),
    .o(al_34c94edb));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_8d03cc1 (
    .a(al_83ae9a40),
    .b(al_6db5b9d2),
    .c(al_4f6bae56[2]),
    .d(al_4f6bae56[3]),
    .e(al_4f6bae56[4]),
    .f(al_4f6bae56[5]),
    .o(al_f60ec0d5));
  AL_DFF_0 al_e6ac790b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9609a6f5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f6bae56[0]));
  AL_DFF_0 al_f9c622ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bf0c650),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f6bae56[1]));
  AL_DFF_0 al_deb482a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f7a09f99),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_206e4ef2[2]));
  AL_DFF_0 al_fc52e269 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_116d91a8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_206e4ef2[3]));
  AL_DFF_0 al_3887fc99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3197cad9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_206e4ef2[4]));
  AL_DFF_0 al_8f6b41a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8f13de6b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_206e4ef2[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_f22c03bb (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_206e4ef2[0]),
    .e(al_206e4ef2[1]),
    .f(al_206e4ef2[2]),
    .o(al_d7967164));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_6bbaec06 (
    .a(al_d7967164),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_206e4ef2[3]),
    .f(al_206e4ef2[4]),
    .o(al_c5c99a19));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_164cadff (
    .a(al_c5c99a19),
    .b(al_206e4ef2[5]),
    .c(al_a48594d3),
    .d(al_4caca369[0]),
    .o(al_dc9abd46));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_9d85af2a (
    .a(al_dc9abd46),
    .b(al_206e4ef2[0]),
    .c(al_206e4ef2[1]),
    .o(al_8f5d07af));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_4e887e50 (
    .a(al_8f5d07af),
    .b(al_6db5b9d2),
    .c(al_206e4ef2[2]),
    .d(al_206e4ef2[3]),
    .e(al_206e4ef2[4]),
    .o(al_3197cad9));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_60c3d3cb (
    .a(al_8f5d07af),
    .b(al_6db5b9d2),
    .c(al_206e4ef2[2]),
    .d(al_206e4ef2[3]),
    .o(al_116d91a8));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_ebfc9d2f (
    .a(al_dc9abd46),
    .b(al_6db5b9d2),
    .c(al_206e4ef2[0]),
    .o(al_56102450));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_45008494 (
    .a(al_dc9abd46),
    .b(al_6db5b9d2),
    .c(al_206e4ef2[0]),
    .d(al_206e4ef2[1]),
    .o(al_ddf07c29));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_c4b129bd (
    .a(al_8f5d07af),
    .b(al_6db5b9d2),
    .c(al_206e4ef2[2]),
    .o(al_f7a09f99));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_67afee58 (
    .a(al_8f5d07af),
    .b(al_6db5b9d2),
    .c(al_206e4ef2[2]),
    .d(al_206e4ef2[3]),
    .e(al_206e4ef2[4]),
    .f(al_206e4ef2[5]),
    .o(al_8f13de6b));
  AL_DFF_0 al_91b76484 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56102450),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_206e4ef2[0]));
  AL_DFF_0 al_625060fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ddf07c29),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_206e4ef2[1]));
  AL_DFF_0 al_4b9e8320 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a7c305cd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ead25ba5[2]));
  AL_DFF_0 al_2b18feb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_32307526),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ead25ba5[3]));
  AL_DFF_0 al_d0a97e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ddc0b8a6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ead25ba5[4]));
  AL_DFF_0 al_bf018e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ab813978),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ead25ba5[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_97e721be (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_ead25ba5[0]),
    .e(al_ead25ba5[1]),
    .f(al_ead25ba5[2]),
    .o(al_c66db911));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_6a0535c8 (
    .a(al_c66db911),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_ead25ba5[3]),
    .f(al_ead25ba5[4]),
    .o(al_2cac5213));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_b3ba110c (
    .a(al_2cac5213),
    .b(al_ead25ba5[5]),
    .c(al_521fd670),
    .d(al_b065182c[0]),
    .o(al_52694b4b));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_eba8896f (
    .a(al_52694b4b),
    .b(al_ead25ba5[0]),
    .c(al_ead25ba5[1]),
    .o(al_bd85c50d));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_5c373186 (
    .a(al_bd85c50d),
    .b(al_6db5b9d2),
    .c(al_ead25ba5[2]),
    .d(al_ead25ba5[3]),
    .e(al_ead25ba5[4]),
    .o(al_ddc0b8a6));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_9b9f7da9 (
    .a(al_bd85c50d),
    .b(al_6db5b9d2),
    .c(al_ead25ba5[2]),
    .d(al_ead25ba5[3]),
    .o(al_32307526));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_15f3d4e (
    .a(al_52694b4b),
    .b(al_6db5b9d2),
    .c(al_ead25ba5[0]),
    .o(al_2a43f573));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_f60c3a39 (
    .a(al_52694b4b),
    .b(al_6db5b9d2),
    .c(al_ead25ba5[0]),
    .d(al_ead25ba5[1]),
    .o(al_9752d581));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_ace637bd (
    .a(al_bd85c50d),
    .b(al_6db5b9d2),
    .c(al_ead25ba5[2]),
    .o(al_a7c305cd));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_6a1b2a15 (
    .a(al_bd85c50d),
    .b(al_6db5b9d2),
    .c(al_ead25ba5[2]),
    .d(al_ead25ba5[3]),
    .e(al_ead25ba5[4]),
    .f(al_ead25ba5[5]),
    .o(al_ab813978));
  AL_DFF_0 al_114545a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2a43f573),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ead25ba5[0]));
  AL_DFF_0 al_cd91993f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9752d581),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ead25ba5[1]));
  AL_DFF_0 al_a8af9eb6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_21a638b3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b04a4cbc[2]));
  AL_DFF_0 al_e9ab30aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3d90e9a3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b04a4cbc[3]));
  AL_DFF_0 al_56a22bab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e377f7a4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b04a4cbc[4]));
  AL_DFF_0 al_8798880b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7cf355db),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b04a4cbc[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_a0316ccd (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_b04a4cbc[0]),
    .e(al_b04a4cbc[1]),
    .f(al_b04a4cbc[2]),
    .o(al_b7e19172));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_a4517ac1 (
    .a(al_b7e19172),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_b04a4cbc[3]),
    .f(al_b04a4cbc[4]),
    .o(al_9e2fe654));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_be95e0a6 (
    .a(al_9e2fe654),
    .b(al_b04a4cbc[5]),
    .c(al_1919cac5),
    .d(al_28515a17[0]),
    .o(al_b6ed5e1b));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_5de20abd (
    .a(al_b6ed5e1b),
    .b(al_b04a4cbc[0]),
    .c(al_b04a4cbc[1]),
    .o(al_63293fc5));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_ebee38eb (
    .a(al_63293fc5),
    .b(al_6db5b9d2),
    .c(al_b04a4cbc[2]),
    .d(al_b04a4cbc[3]),
    .e(al_b04a4cbc[4]),
    .o(al_e377f7a4));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_3d0bb20a (
    .a(al_63293fc5),
    .b(al_6db5b9d2),
    .c(al_b04a4cbc[2]),
    .d(al_b04a4cbc[3]),
    .o(al_3d90e9a3));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_4ba66268 (
    .a(al_b6ed5e1b),
    .b(al_6db5b9d2),
    .c(al_b04a4cbc[0]),
    .o(al_13f5c59d));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_b04c80ca (
    .a(al_b6ed5e1b),
    .b(al_6db5b9d2),
    .c(al_b04a4cbc[0]),
    .d(al_b04a4cbc[1]),
    .o(al_7329b916));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_3669efed (
    .a(al_63293fc5),
    .b(al_6db5b9d2),
    .c(al_b04a4cbc[2]),
    .o(al_21a638b3));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_a13533a8 (
    .a(al_63293fc5),
    .b(al_6db5b9d2),
    .c(al_b04a4cbc[2]),
    .d(al_b04a4cbc[3]),
    .e(al_b04a4cbc[4]),
    .f(al_b04a4cbc[5]),
    .o(al_7cf355db));
  AL_DFF_0 al_b545fc09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_13f5c59d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b04a4cbc[0]));
  AL_DFF_0 al_853f7609 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7329b916),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b04a4cbc[1]));
  AL_DFF_0 al_4909a7af (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ec64ca16),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b9e1d84[2]));
  AL_DFF_0 al_5580bad4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ebf34b40),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b9e1d84[3]));
  AL_DFF_0 al_e7a255ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aeeedc7e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b9e1d84[4]));
  AL_DFF_0 al_74e468b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_42eb8568),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b9e1d84[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_6f03d87a (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_6b9e1d84[0]),
    .e(al_6b9e1d84[1]),
    .f(al_6b9e1d84[2]),
    .o(al_7ab8db7c));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_1ee06792 (
    .a(al_7ab8db7c),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_6b9e1d84[3]),
    .f(al_6b9e1d84[4]),
    .o(al_be012e15));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_10d36531 (
    .a(al_be012e15),
    .b(al_6b9e1d84[5]),
    .c(al_6e50ac65),
    .d(al_28515a17[0]),
    .o(al_8ec0a0c8));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_af037b9e (
    .a(al_8ec0a0c8),
    .b(al_6b9e1d84[0]),
    .c(al_6b9e1d84[1]),
    .d(al_6b9e1d84[2]),
    .e(al_6b9e1d84[3]),
    .f(al_6b9e1d84[4]),
    .o(al_acd1c245));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_1857da1f (
    .a(al_8ec0a0c8),
    .b(al_6b9e1d84[0]),
    .c(al_6b9e1d84[1]),
    .d(al_6b9e1d84[2]),
    .e(al_6b9e1d84[3]),
    .f(al_6b9e1d84[4]),
    .o(al_5477c30f));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_f6601305 (
    .a(al_5477c30f),
    .b(al_6db5b9d2),
    .o(al_aeeedc7e));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_76ae900b (
    .a(al_8ec0a0c8),
    .b(al_6db5b9d2),
    .c(al_6b9e1d84[0]),
    .d(al_6b9e1d84[1]),
    .e(al_6b9e1d84[2]),
    .f(al_6b9e1d84[3]),
    .o(al_ebf34b40));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_742b0374 (
    .a(al_8ec0a0c8),
    .b(al_6db5b9d2),
    .c(al_6b9e1d84[0]),
    .o(al_aff4e477));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_6e79ed7f (
    .a(al_8ec0a0c8),
    .b(al_6db5b9d2),
    .c(al_6b9e1d84[0]),
    .d(al_6b9e1d84[1]),
    .o(al_e7777d0d));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_3b75396b (
    .a(al_8ec0a0c8),
    .b(al_6db5b9d2),
    .c(al_6b9e1d84[0]),
    .d(al_6b9e1d84[1]),
    .e(al_6b9e1d84[2]),
    .o(al_ec64ca16));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_c66b2f15 (
    .a(al_acd1c245),
    .b(al_6db5b9d2),
    .c(al_6b9e1d84[5]),
    .o(al_42eb8568));
  AL_DFF_0 al_34e1eb76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aff4e477),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b9e1d84[0]));
  AL_DFF_0 al_af578eed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e7777d0d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b9e1d84[1]));
  AL_DFF_0 al_e0d9a5f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_61e4c12),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c244bf8b[2]));
  AL_DFF_0 al_ffebafe1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e75ba485),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c244bf8b[3]));
  AL_DFF_0 al_4e2216b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_594d9eef),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c244bf8b[4]));
  AL_DFF_0 al_86a03e60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f6290e5d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c244bf8b[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_8b4e0fb0 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_c244bf8b[0]),
    .e(al_c244bf8b[1]),
    .f(al_c244bf8b[2]),
    .o(al_994a49f));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_c6c194a7 (
    .a(al_994a49f),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_c244bf8b[3]),
    .f(al_c244bf8b[4]),
    .o(al_957b61e0));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_5665626b (
    .a(al_957b61e0),
    .b(al_c244bf8b[5]),
    .c(al_8dc56974),
    .d(al_4caca369[0]),
    .o(al_9f34fb19));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_61c56357 (
    .a(al_9f34fb19),
    .b(al_c244bf8b[0]),
    .c(al_c244bf8b[1]),
    .o(al_e96a29f2));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_6d61180d (
    .a(al_e96a29f2),
    .b(al_6db5b9d2),
    .c(al_c244bf8b[2]),
    .d(al_c244bf8b[3]),
    .e(al_c244bf8b[4]),
    .o(al_594d9eef));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_3b92468b (
    .a(al_e96a29f2),
    .b(al_6db5b9d2),
    .c(al_c244bf8b[2]),
    .d(al_c244bf8b[3]),
    .o(al_e75ba485));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_5a404b8a (
    .a(al_9f34fb19),
    .b(al_6db5b9d2),
    .c(al_c244bf8b[0]),
    .o(al_fd1d15be));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_b6ab7e43 (
    .a(al_9f34fb19),
    .b(al_6db5b9d2),
    .c(al_c244bf8b[0]),
    .d(al_c244bf8b[1]),
    .o(al_7f125c63));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_3ab611f6 (
    .a(al_e96a29f2),
    .b(al_6db5b9d2),
    .c(al_c244bf8b[2]),
    .o(al_61e4c12));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_a7f0123e (
    .a(al_e96a29f2),
    .b(al_6db5b9d2),
    .c(al_c244bf8b[2]),
    .d(al_c244bf8b[3]),
    .e(al_c244bf8b[4]),
    .f(al_c244bf8b[5]),
    .o(al_f6290e5d));
  AL_DFF_0 al_72e95d42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fd1d15be),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c244bf8b[0]));
  AL_DFF_0 al_7508efd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7f125c63),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c244bf8b[1]));
  AL_DFF_0 al_7047c74f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_27647c5b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d44a73a0[2]));
  AL_DFF_0 al_856953a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_359de7f7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d44a73a0[3]));
  AL_DFF_0 al_74532b39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_84cbc97b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d44a73a0[4]));
  AL_DFF_0 al_f7eb6e61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a2e27860),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d44a73a0[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_f4adf795 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_d44a73a0[0]),
    .e(al_d44a73a0[1]),
    .f(al_d44a73a0[2]),
    .o(al_65ea04b6));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_8f9d9160 (
    .a(al_65ea04b6),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_d44a73a0[3]),
    .f(al_d44a73a0[4]),
    .o(al_ba6805c2));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_512a3f62 (
    .a(al_ba6805c2),
    .b(al_d44a73a0[5]),
    .c(al_8b05cae6),
    .d(al_b065182c[0]),
    .o(al_29e29c2));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_59dd1534 (
    .a(al_29e29c2),
    .b(al_d44a73a0[0]),
    .c(al_d44a73a0[1]),
    .o(al_3fb2454f));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_f3ebbb9e (
    .a(al_3fb2454f),
    .b(al_6db5b9d2),
    .c(al_d44a73a0[2]),
    .d(al_d44a73a0[3]),
    .e(al_d44a73a0[4]),
    .o(al_84cbc97b));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_7f05c302 (
    .a(al_3fb2454f),
    .b(al_6db5b9d2),
    .c(al_d44a73a0[2]),
    .d(al_d44a73a0[3]),
    .o(al_359de7f7));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_974b8788 (
    .a(al_29e29c2),
    .b(al_6db5b9d2),
    .c(al_d44a73a0[0]),
    .o(al_e0bee367));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_1f5416b4 (
    .a(al_29e29c2),
    .b(al_6db5b9d2),
    .c(al_d44a73a0[0]),
    .d(al_d44a73a0[1]),
    .o(al_ad44d351));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_8a2381a (
    .a(al_3fb2454f),
    .b(al_6db5b9d2),
    .c(al_d44a73a0[2]),
    .o(al_27647c5b));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_90a29ca3 (
    .a(al_3fb2454f),
    .b(al_6db5b9d2),
    .c(al_d44a73a0[2]),
    .d(al_d44a73a0[3]),
    .e(al_d44a73a0[4]),
    .f(al_d44a73a0[5]),
    .o(al_a2e27860));
  AL_DFF_0 al_ccd76124 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e0bee367),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d44a73a0[0]));
  AL_DFF_0 al_d38ac002 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ad44d351),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d44a73a0[1]));
  AL_DFF_0 al_ef385a29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bc75ce6f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_37663fe4[2]));
  AL_DFF_0 al_5cb9878a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4a9b23a9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_37663fe4[3]));
  AL_DFF_0 al_39019cde (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cee52ae5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_37663fe4[4]));
  AL_DFF_0 al_2c76dad4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ad9326a7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_37663fe4[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_364ac2c8 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_37663fe4[0]),
    .e(al_37663fe4[1]),
    .f(al_37663fe4[2]),
    .o(al_4743910a));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_6366d9d (
    .a(al_4743910a),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_37663fe4[3]),
    .f(al_37663fe4[4]),
    .o(al_7905d584));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_dfeea24f (
    .a(al_7905d584),
    .b(al_37663fe4[5]),
    .c(al_7bafa36d),
    .d(al_28515a17[0]),
    .o(al_3c305c5d));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_c077a722 (
    .a(al_3c305c5d),
    .b(al_37663fe4[0]),
    .c(al_37663fe4[1]),
    .o(al_d77438af));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_b6a10136 (
    .a(al_d77438af),
    .b(al_6db5b9d2),
    .c(al_37663fe4[2]),
    .d(al_37663fe4[3]),
    .e(al_37663fe4[4]),
    .o(al_cee52ae5));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_d26259d8 (
    .a(al_d77438af),
    .b(al_6db5b9d2),
    .c(al_37663fe4[2]),
    .d(al_37663fe4[3]),
    .o(al_4a9b23a9));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_9b0746bf (
    .a(al_3c305c5d),
    .b(al_6db5b9d2),
    .c(al_37663fe4[0]),
    .o(al_47d4f942));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_3ef859f7 (
    .a(al_3c305c5d),
    .b(al_6db5b9d2),
    .c(al_37663fe4[0]),
    .d(al_37663fe4[1]),
    .o(al_b7074965));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_99898e16 (
    .a(al_d77438af),
    .b(al_6db5b9d2),
    .c(al_37663fe4[2]),
    .o(al_bc75ce6f));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_8fb8f328 (
    .a(al_d77438af),
    .b(al_6db5b9d2),
    .c(al_37663fe4[2]),
    .d(al_37663fe4[3]),
    .e(al_37663fe4[4]),
    .f(al_37663fe4[5]),
    .o(al_ad9326a7));
  AL_DFF_0 al_66c26ab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_47d4f942),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_37663fe4[0]));
  AL_DFF_0 al_c12ddbe9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7074965),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_37663fe4[1]));
  AL_DFF_0 al_9e2b0728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b04b1b3b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[0]));
  AL_DFF_0 al_9e79b36b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b04b1b3b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[1]));
  AL_DFF_0 al_21e5a258 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b04b1b3b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[2]));
  AL_DFF_0 al_3cc943c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b04b1b3b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[3]));
  AL_DFF_0 al_487928d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b04b1b3b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[4]));
  AL_DFF_0 al_689ed924 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b04b1b3b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[5]));
  AL_DFF_0 al_b2f9c52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea67686c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[6]));
  AL_DFF_0 al_2ca0e080 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea67686c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[7]));
  AL_DFF_0 al_c337cefe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea67686c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[8]));
  AL_DFF_0 al_58a2a317 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea67686c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[9]));
  AL_DFF_0 al_f4d09cce (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea67686c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[10]));
  AL_DFF_0 al_d62727fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea67686c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[11]));
  AL_DFF_0 al_bf773934 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_27ec7185[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[12]));
  AL_DFF_0 al_153ab70c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_27ec7185[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[13]));
  AL_DFF_0 al_e7e2e941 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_27ec7185[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[14]));
  AL_DFF_0 al_ae558272 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_27ec7185[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[15]));
  AL_DFF_0 al_89bfd912 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_27ec7185[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[16]));
  AL_DFF_0 al_4efaf1d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_27ec7185[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[17]));
  AL_DFF_0 al_ccc417ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5342096[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[18]));
  AL_DFF_0 al_3588f57d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5342096[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[19]));
  AL_DFF_0 al_d479565f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5342096[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[20]));
  AL_DFF_0 al_68627895 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5342096[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[21]));
  AL_DFF_0 al_28aee54b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5342096[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[22]));
  AL_DFF_0 al_5f46a73b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5342096[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[23]));
  AL_DFF_0 al_293fe346 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a84549[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[24]));
  AL_DFF_0 al_aad3c098 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a84549[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[25]));
  AL_DFF_0 al_9b3df5ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a84549[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[26]));
  AL_DFF_0 al_1b0a0585 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a84549[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[27]));
  AL_DFF_0 al_26a6fe12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a84549[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[28]));
  AL_DFF_0 al_16c723d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5a84549[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[29]));
  AL_DFF_0 al_f379ecab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_764d3602[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[30]));
  AL_DFF_0 al_69f92934 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_764d3602[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[31]));
  AL_DFF_0 al_2445e3d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_764d3602[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[32]));
  AL_DFF_0 al_88c13fdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_764d3602[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[33]));
  AL_DFF_0 al_af8eaa93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_764d3602[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[34]));
  AL_DFF_0 al_3d0f4d74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_764d3602[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[35]));
  AL_DFF_0 al_1f1a5624 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9bc4f0be[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[36]));
  AL_DFF_0 al_521ad6f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9bc4f0be[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[37]));
  AL_DFF_0 al_8348e98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9bc4f0be[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[38]));
  AL_DFF_0 al_465477a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9bc4f0be[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[39]));
  AL_DFF_0 al_2efab1d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9bc4f0be[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[40]));
  AL_DFF_0 al_fb927ffd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9bc4f0be[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[41]));
  AL_DFF_0 al_ca23b3a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9427b946[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[42]));
  AL_DFF_0 al_33a74fbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9427b946[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[43]));
  AL_DFF_0 al_5b0b6694 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9427b946[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[44]));
  AL_DFF_0 al_896ffa9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9427b946[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[45]));
  AL_DFF_0 al_7d1952e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9427b946[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[46]));
  AL_DFF_0 al_546a5c1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9427b946[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[47]));
  AL_DFF_0 al_eb3fec6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6a612a6[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[48]));
  AL_DFF_0 al_83e7b746 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6a612a6[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[49]));
  AL_DFF_0 al_72d62682 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6a612a6[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[50]));
  AL_DFF_0 al_2bf5f308 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6a612a6[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[51]));
  AL_DFF_0 al_34c20063 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6a612a6[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[52]));
  AL_DFF_0 al_8558a088 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6a612a6[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[53]));
  AL_DFF_0 al_8b4bba41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_92e7eeea[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[54]));
  AL_DFF_0 al_6a0823bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_92e7eeea[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[55]));
  AL_DFF_0 al_245b4066 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_92e7eeea[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[56]));
  AL_DFF_0 al_ff6102c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_92e7eeea[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[57]));
  AL_DFF_0 al_ab56b6ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_92e7eeea[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[58]));
  AL_DFF_0 al_d631a522 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_92e7eeea[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[59]));
  AL_DFF_0 al_667233f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b48e0e9a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[60]));
  AL_DFF_0 al_53453e1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b48e0e9a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[61]));
  AL_DFF_0 al_d90e9fe1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b48e0e9a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[62]));
  AL_DFF_0 al_14c50921 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b48e0e9a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[63]));
  AL_DFF_0 al_81a49484 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b48e0e9a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[64]));
  AL_DFF_0 al_d60a5ed4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b48e0e9a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[65]));
  AL_DFF_0 al_65ca24dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_175c7e02[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[66]));
  AL_DFF_0 al_908f9edb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_175c7e02[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[67]));
  AL_DFF_0 al_5e63bf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_175c7e02[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[68]));
  AL_DFF_0 al_4019debf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_175c7e02[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[69]));
  AL_DFF_0 al_a4c9857e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_175c7e02[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[70]));
  AL_DFF_0 al_f0b8961 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_175c7e02[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[71]));
  AL_DFF_0 al_affcaf9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33614149[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[72]));
  AL_DFF_0 al_64dc3fda (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33614149[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[73]));
  AL_DFF_0 al_3d783422 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33614149[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[74]));
  AL_DFF_0 al_a1d3c01e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33614149[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[75]));
  AL_DFF_0 al_dfc54cf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33614149[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[76]));
  AL_DFF_0 al_36f0c9a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33614149[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[77]));
  AL_DFF_0 al_3427d1c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ed19afe1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[78]));
  AL_DFF_0 al_7321112e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ed19afe1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[79]));
  AL_DFF_0 al_b20d2262 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ed19afe1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[80]));
  AL_DFF_0 al_61b90edb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ed19afe1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[81]));
  AL_DFF_0 al_7454058b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ed19afe1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[82]));
  AL_DFF_0 al_1fdd2bbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ed19afe1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[83]));
  AL_DFF_0 al_3e6a2383 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_87305132[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[84]));
  AL_DFF_0 al_f8b79d1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_87305132[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[85]));
  AL_DFF_0 al_f4257cf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_87305132[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[86]));
  AL_DFF_0 al_cc118c33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_87305132[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[87]));
  AL_DFF_0 al_cd4d90ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_87305132[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[88]));
  AL_DFF_0 al_70ea54a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_87305132[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[89]));
  AL_DFF_0 al_b15e5d55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fce7b5a9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[90]));
  AL_DFF_0 al_bf721059 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fce7b5a9[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[91]));
  AL_DFF_0 al_d1e73e99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fce7b5a9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[92]));
  AL_DFF_0 al_305dbf69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fce7b5a9[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[93]));
  AL_DFF_0 al_bc374fea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fce7b5a9[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[94]));
  AL_DFF_0 al_7a029a0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fce7b5a9[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[95]));
  AL_DFF_0 al_38f1f7e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_407652d9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[96]));
  AL_DFF_0 al_5e36e663 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_407652d9[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[97]));
  AL_DFF_0 al_8556888e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_407652d9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[98]));
  AL_DFF_0 al_ebee031a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_407652d9[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[99]));
  AL_DFF_0 al_cc507c62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_407652d9[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[100]));
  AL_DFF_0 al_2a06f000 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_407652d9[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[101]));
  AL_DFF_0 al_6fe843d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c527aa4e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[102]));
  AL_DFF_0 al_5508d834 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c527aa4e[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[103]));
  AL_DFF_0 al_a2a5c915 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c527aa4e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[104]));
  AL_DFF_0 al_feab3af3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c527aa4e[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[105]));
  AL_DFF_0 al_d9e1e5e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c527aa4e[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[106]));
  AL_DFF_0 al_7e42536 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c527aa4e[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[107]));
  AL_DFF_0 al_dae03da1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7a189[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[108]));
  AL_DFF_0 al_978e98f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7a189[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[109]));
  AL_DFF_0 al_3c0503b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7a189[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[110]));
  AL_DFF_0 al_124d5e8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7a189[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[111]));
  AL_DFF_0 al_2af70e3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7a189[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[112]));
  AL_DFF_0 al_1dacfda7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7a189[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[113]));
  AL_DFF_0 al_b3f4428 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_63020263[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[114]));
  AL_DFF_0 al_f2d6fa22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_63020263[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[115]));
  AL_DFF_0 al_742e9905 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_63020263[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[116]));
  AL_DFF_0 al_dd3c8777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_63020263[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[117]));
  AL_DFF_0 al_b023653f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_63020263[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[118]));
  AL_DFF_0 al_81121501 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_63020263[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[119]));
  AL_DFF_0 al_a7698580 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98058573[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[120]));
  AL_DFF_0 al_f0f32d18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98058573[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[121]));
  AL_DFF_0 al_6277fa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98058573[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[122]));
  AL_DFF_0 al_336f29b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98058573[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[123]));
  AL_DFF_0 al_ca74cb41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98058573[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[124]));
  AL_DFF_0 al_8abd65c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98058573[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[125]));
  AL_DFF_0 al_84dba6c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69204309[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[126]));
  AL_DFF_0 al_94f19d96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69204309[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[127]));
  AL_DFF_0 al_b0096c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69204309[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[128]));
  AL_DFF_0 al_2a435981 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69204309[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[129]));
  AL_DFF_0 al_bdd1c253 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69204309[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[130]));
  AL_DFF_0 al_85f15dbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69204309[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[131]));
  AL_DFF_0 al_1b39c26c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9ca6681[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[132]));
  AL_DFF_0 al_901c1109 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9ca6681[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[133]));
  AL_DFF_0 al_b2222d09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9ca6681[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[134]));
  AL_DFF_0 al_7675f901 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9ca6681[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[135]));
  AL_DFF_0 al_d3ef48e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9ca6681[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[136]));
  AL_DFF_0 al_aca1967f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9ca6681[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[137]));
  AL_DFF_0 al_ede57b75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a5ad4b3c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[138]));
  AL_DFF_0 al_3a8964ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a5ad4b3c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[139]));
  AL_DFF_0 al_b2d46147 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a5ad4b3c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[140]));
  AL_DFF_0 al_6dd5b513 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a5ad4b3c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[141]));
  AL_DFF_0 al_7d1116b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a5ad4b3c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[142]));
  AL_DFF_0 al_3fac87d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a5ad4b3c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[143]));
  AL_DFF_0 al_15141922 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3a9b666[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[144]));
  AL_DFF_0 al_32f663df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3a9b666[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[145]));
  AL_DFF_0 al_fa5224d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3a9b666[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[146]));
  AL_DFF_0 al_fca1da2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3a9b666[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[147]));
  AL_DFF_0 al_84e3ffb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3a9b666[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[148]));
  AL_DFF_0 al_f31a7589 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3a9b666[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[149]));
  AL_DFF_0 al_d09af4bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f033fc44[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[150]));
  AL_DFF_0 al_b5fe9665 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f033fc44[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[151]));
  AL_DFF_0 al_d9918c13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f033fc44[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[152]));
  AL_DFF_0 al_a2095087 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f033fc44[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[153]));
  AL_DFF_0 al_9ba280c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f033fc44[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[154]));
  AL_DFF_0 al_3ee25ad8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f033fc44[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[155]));
  AL_DFF_0 al_fccc0f75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b8da42f7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[156]));
  AL_DFF_0 al_e3f7cffc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b8da42f7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[157]));
  AL_DFF_0 al_3fc09254 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b8da42f7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[158]));
  AL_DFF_0 al_c1bbc455 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b8da42f7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[159]));
  AL_DFF_0 al_afd9d801 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b8da42f7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[160]));
  AL_DFF_0 al_5747d59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b8da42f7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[161]));
  AL_DFF_0 al_30af378a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d88fcc0f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[162]));
  AL_DFF_0 al_3abe1832 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d88fcc0f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[163]));
  AL_DFF_0 al_3e06e0bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d88fcc0f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[164]));
  AL_DFF_0 al_375e487 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d88fcc0f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[165]));
  AL_DFF_0 al_29066105 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d88fcc0f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[166]));
  AL_DFF_0 al_ba699ea4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d88fcc0f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[167]));
  AL_DFF_0 al_fb79f68b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b88a45c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[168]));
  AL_DFF_0 al_d8d3475a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b88a45c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[169]));
  AL_DFF_0 al_7bdc57a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b88a45c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[170]));
  AL_DFF_0 al_b0db64d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b88a45c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[171]));
  AL_DFF_0 al_fc627b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b88a45c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[172]));
  AL_DFF_0 al_74e714bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8b88a45c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[173]));
  AL_DFF_0 al_aa741f26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c25a985[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[174]));
  AL_DFF_0 al_a7270c9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c25a985[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[175]));
  AL_DFF_0 al_523f956b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c25a985[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[176]));
  AL_DFF_0 al_b2d34ecd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c25a985[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[177]));
  AL_DFF_0 al_1265a314 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c25a985[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[178]));
  AL_DFF_0 al_b1a924cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c25a985[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[179]));
  AL_DFF_0 al_74018ad9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2c2ca002[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[180]));
  AL_DFF_0 al_1b617045 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2c2ca002[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[181]));
  AL_DFF_0 al_5ef9f601 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2c2ca002[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[182]));
  AL_DFF_0 al_d54a339d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2c2ca002[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[183]));
  AL_DFF_0 al_c29b2a83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2c2ca002[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[184]));
  AL_DFF_0 al_a01133e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2c2ca002[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[185]));
  AL_DFF_0 al_b631655e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d0d403d6[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[186]));
  AL_DFF_0 al_d15b6592 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d0d403d6[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[187]));
  AL_DFF_0 al_1a6b948b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d0d403d6[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[188]));
  AL_DFF_0 al_938997cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d0d403d6[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[189]));
  AL_DFF_0 al_c6a02855 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d0d403d6[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[190]));
  AL_DFF_0 al_ab20214e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d0d403d6[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[191]));
  AL_DFF_0 al_e5097e08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3aa16a9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[192]));
  AL_DFF_0 al_e5a4136e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3aa16a9[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[193]));
  AL_DFF_0 al_1000e7fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3aa16a9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[194]));
  AL_DFF_0 al_a8f48204 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3aa16a9[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[195]));
  AL_DFF_0 al_90c2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3aa16a9[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[196]));
  AL_DFF_0 al_96f3aa8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3aa16a9[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[197]));
  AL_DFF_0 al_a5b651a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c1bada4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[198]));
  AL_DFF_0 al_b52ccbd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c1bada4[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[199]));
  AL_DFF_0 al_cbce3922 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c1bada4[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[200]));
  AL_DFF_0 al_2b0d6b0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c1bada4[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[201]));
  AL_DFF_0 al_a7d87f66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c1bada4[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[202]));
  AL_DFF_0 al_117e5d02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4c1bada4[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[203]));
  AL_DFF_0 al_8a582b82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6b6ef69[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[204]));
  AL_DFF_0 al_6b0589fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6b6ef69[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[205]));
  AL_DFF_0 al_420f8d99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6b6ef69[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[206]));
  AL_DFF_0 al_83f36607 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6b6ef69[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[207]));
  AL_DFF_0 al_ff0a6b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6b6ef69[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[208]));
  AL_DFF_0 al_645db5a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6b6ef69[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[209]));
  AL_DFF_0 al_f2ebc1ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0408eb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[210]));
  AL_DFF_0 al_2ef53bae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0408eb[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[211]));
  AL_DFF_0 al_f4e38aa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0408eb[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[212]));
  AL_DFF_0 al_fb4fe877 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0408eb[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[213]));
  AL_DFF_0 al_d2ccd62d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0408eb[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[214]));
  AL_DFF_0 al_d04f1f9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b0408eb[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[215]));
  AL_DFF_0 al_13ff570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5577a41[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[216]));
  AL_DFF_0 al_225fc6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5577a41[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[217]));
  AL_DFF_0 al_856aa183 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5577a41[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[218]));
  AL_DFF_0 al_1710635e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5577a41[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[219]));
  AL_DFF_0 al_1085911 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5577a41[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[220]));
  AL_DFF_0 al_2898e4c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5577a41[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[221]));
  AL_DFF_0 al_eac5be65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d55b2543[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[222]));
  AL_DFF_0 al_431496d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d55b2543[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[223]));
  AL_DFF_0 al_680d177d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d55b2543[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[224]));
  AL_DFF_0 al_851f7cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d55b2543[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[225]));
  AL_DFF_0 al_aa6b5f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d55b2543[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[226]));
  AL_DFF_0 al_d831ba9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d55b2543[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[227]));
  AL_DFF_0 al_5c87acf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0d076bb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[228]));
  AL_DFF_0 al_f9dba3d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0d076bb[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[229]));
  AL_DFF_0 al_f368afac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0d076bb[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[230]));
  AL_DFF_0 al_ead2a302 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0d076bb[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[231]));
  AL_DFF_0 al_67409011 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0d076bb[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[232]));
  AL_DFF_0 al_1bcb4703 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c0d076bb[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[233]));
  AL_DFF_0 al_3767bb9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98c6a23b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[234]));
  AL_DFF_0 al_df67b35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98c6a23b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[235]));
  AL_DFF_0 al_6be41185 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98c6a23b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[236]));
  AL_DFF_0 al_b90f064a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98c6a23b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[237]));
  AL_DFF_0 al_7247e86a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98c6a23b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[238]));
  AL_DFF_0 al_73a7474d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98c6a23b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[239]));
  AL_DFF_0 al_598412b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_77d19440[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[240]));
  AL_DFF_0 al_746969c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_77d19440[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[241]));
  AL_DFF_0 al_82e8a102 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_77d19440[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[242]));
  AL_DFF_0 al_e20873c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_77d19440[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[243]));
  AL_DFF_0 al_80ca1d15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_77d19440[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[244]));
  AL_DFF_0 al_1effeab8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_77d19440[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[245]));
  AL_DFF_0 al_8b47a25b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3fa002d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[246]));
  AL_DFF_0 al_f6f0c9f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3fa002d[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[247]));
  AL_DFF_0 al_de8fc338 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3fa002d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[248]));
  AL_DFF_0 al_580d14c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3fa002d[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[249]));
  AL_DFF_0 al_e01841c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3fa002d[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[250]));
  AL_DFF_0 al_f7d7dfe5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3fa002d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[251]));
  AL_DFF_0 al_c8eee9c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3ab36424[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[252]));
  AL_DFF_0 al_b0005744 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3ab36424[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[253]));
  AL_DFF_0 al_23ad5c22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3ab36424[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[254]));
  AL_DFF_0 al_12dfbd11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3ab36424[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(ddr_app_rd_data[255]));
  AL_DFF_0 al_850c4962 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4cb51ed9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e865b87a[2]));
  AL_DFF_0 al_4e334e31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_efc69db4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e865b87a[3]));
  AL_DFF_0 al_31a500c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_969bce5a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e865b87a[4]));
  AL_DFF_0 al_e4eded5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5bb4cdbf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e865b87a[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_a737e337 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_e865b87a[0]),
    .e(al_e865b87a[1]),
    .f(al_e865b87a[2]),
    .o(al_4fcbf6ef));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_eb6d8b44 (
    .a(al_4fcbf6ef),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_e865b87a[3]),
    .f(al_e865b87a[4]),
    .o(al_b62a0a78));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_18c7adef (
    .a(al_b62a0a78),
    .b(al_e865b87a[5]),
    .c(al_25e4ab96),
    .d(al_4caca369[0]),
    .o(al_466952a1));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_9e7920c1 (
    .a(al_466952a1),
    .b(al_e865b87a[0]),
    .c(al_e865b87a[1]),
    .o(al_6e5cc87d));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_f9ab6e98 (
    .a(al_6e5cc87d),
    .b(al_6db5b9d2),
    .c(al_e865b87a[2]),
    .d(al_e865b87a[3]),
    .e(al_e865b87a[4]),
    .o(al_969bce5a));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_9af5e305 (
    .a(al_6e5cc87d),
    .b(al_6db5b9d2),
    .c(al_e865b87a[2]),
    .d(al_e865b87a[3]),
    .o(al_efc69db4));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_e439d39a (
    .a(al_466952a1),
    .b(al_6db5b9d2),
    .c(al_e865b87a[0]),
    .o(al_75ba7c3a));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_c36b7b8d (
    .a(al_466952a1),
    .b(al_6db5b9d2),
    .c(al_e865b87a[0]),
    .d(al_e865b87a[1]),
    .o(al_cf7de8fd));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_824e3da4 (
    .a(al_6e5cc87d),
    .b(al_6db5b9d2),
    .c(al_e865b87a[2]),
    .o(al_4cb51ed9));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_7404a5d3 (
    .a(al_6e5cc87d),
    .b(al_6db5b9d2),
    .c(al_e865b87a[2]),
    .d(al_e865b87a[3]),
    .e(al_e865b87a[4]),
    .f(al_e865b87a[5]),
    .o(al_5bb4cdbf));
  AL_DFF_0 al_f3936f92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_75ba7c3a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e865b87a[0]));
  AL_DFF_0 al_8392fba5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf7de8fd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e865b87a[1]));
  AL_DFF_0 al_d75c19c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_23ffeaf6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f359f0c8[2]));
  AL_DFF_0 al_e71cf3e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ab1a88b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f359f0c8[3]));
  AL_DFF_0 al_f10750b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7ba8863),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f359f0c8[4]));
  AL_DFF_0 al_8f77653 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6a0564ce),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f359f0c8[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_b7a96c (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_f359f0c8[0]),
    .e(al_f359f0c8[1]),
    .f(al_f359f0c8[2]),
    .o(al_ddc5d17a));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_591d1174 (
    .a(al_ddc5d17a),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_f359f0c8[3]),
    .f(al_f359f0c8[4]),
    .o(al_b09bcab2));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_f0bbab71 (
    .a(al_b09bcab2),
    .b(al_f359f0c8[5]),
    .c(al_6e370c03),
    .d(al_b065182c[0]),
    .o(al_e8b6474b));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_b9bcb80a (
    .a(al_e8b6474b),
    .b(al_f359f0c8[0]),
    .c(al_f359f0c8[1]),
    .o(al_f2a9e54d));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_4f47550 (
    .a(al_f2a9e54d),
    .b(al_6db5b9d2),
    .c(al_f359f0c8[2]),
    .d(al_f359f0c8[3]),
    .e(al_f359f0c8[4]),
    .o(al_b7ba8863));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_9d9262c (
    .a(al_f2a9e54d),
    .b(al_6db5b9d2),
    .c(al_f359f0c8[2]),
    .d(al_f359f0c8[3]),
    .o(al_ab1a88b1));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_cf19853c (
    .a(al_e8b6474b),
    .b(al_6db5b9d2),
    .c(al_f359f0c8[0]),
    .o(al_ce51fefb));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_6c3b50a1 (
    .a(al_e8b6474b),
    .b(al_6db5b9d2),
    .c(al_f359f0c8[0]),
    .d(al_f359f0c8[1]),
    .o(al_875002d2));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_c891f154 (
    .a(al_f2a9e54d),
    .b(al_6db5b9d2),
    .c(al_f359f0c8[2]),
    .o(al_23ffeaf6));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_c2001289 (
    .a(al_f2a9e54d),
    .b(al_6db5b9d2),
    .c(al_f359f0c8[2]),
    .d(al_f359f0c8[3]),
    .e(al_f359f0c8[4]),
    .f(al_f359f0c8[5]),
    .o(al_6a0564ce));
  AL_DFF_0 al_e5244e45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ce51fefb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f359f0c8[0]));
  AL_DFF_0 al_3571de60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_875002d2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f359f0c8[1]));
  AL_DFF_0 al_1b16af00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55d82b12),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a14e36[2]));
  AL_DFF_0 al_5bd72066 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_65273b79),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a14e36[3]));
  AL_DFF_0 al_1889afbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_199366db),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a14e36[4]));
  AL_DFF_0 al_1c5319d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e1e03eb2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a14e36[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_ff91a8e9 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_85a14e36[0]),
    .e(al_85a14e36[1]),
    .f(al_85a14e36[2]),
    .o(al_2bfd730a));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_42ca63b5 (
    .a(al_2bfd730a),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_85a14e36[3]),
    .f(al_85a14e36[4]),
    .o(al_c21b49ee));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_ac297d14 (
    .a(al_c21b49ee),
    .b(al_85a14e36[5]),
    .c(al_770f9dd1),
    .d(al_28515a17[0]),
    .o(al_7581b68c));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_d9074990 (
    .a(al_7581b68c),
    .b(al_85a14e36[0]),
    .c(al_85a14e36[1]),
    .o(al_e53fc54d));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_5d4c7dbe (
    .a(al_e53fc54d),
    .b(al_6db5b9d2),
    .c(al_85a14e36[2]),
    .d(al_85a14e36[3]),
    .e(al_85a14e36[4]),
    .o(al_199366db));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_7f7650be (
    .a(al_e53fc54d),
    .b(al_6db5b9d2),
    .c(al_85a14e36[2]),
    .d(al_85a14e36[3]),
    .o(al_65273b79));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_6be2bf84 (
    .a(al_7581b68c),
    .b(al_6db5b9d2),
    .c(al_85a14e36[0]),
    .o(al_36fbd71d));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_18cbc121 (
    .a(al_7581b68c),
    .b(al_6db5b9d2),
    .c(al_85a14e36[0]),
    .d(al_85a14e36[1]),
    .o(al_800e1ab8));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_fec941ef (
    .a(al_e53fc54d),
    .b(al_6db5b9d2),
    .c(al_85a14e36[2]),
    .o(al_55d82b12));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_29c77131 (
    .a(al_e53fc54d),
    .b(al_6db5b9d2),
    .c(al_85a14e36[2]),
    .d(al_85a14e36[3]),
    .e(al_85a14e36[4]),
    .f(al_85a14e36[5]),
    .o(al_e1e03eb2));
  AL_DFF_0 al_5d2abd80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_36fbd71d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a14e36[0]));
  AL_DFF_0 al_e3552960 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_800e1ab8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a14e36[1]));
  AL_DFF_0 al_89a4d2b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_552a02c8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e31889d8[2]));
  AL_DFF_0 al_587592d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_45ef6b15),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e31889d8[3]));
  AL_DFF_0 al_41cf112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_322f98e5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e31889d8[4]));
  AL_DFF_0 al_e28c466 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2684592f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e31889d8[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_ca29925e (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_e31889d8[0]),
    .e(al_e31889d8[1]),
    .f(al_e31889d8[2]),
    .o(al_39c9e6e2));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_b77f4fe8 (
    .a(al_39c9e6e2),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_e31889d8[3]),
    .f(al_e31889d8[4]),
    .o(al_a6be8738));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_82f97a31 (
    .a(al_a6be8738),
    .b(al_e31889d8[5]),
    .c(al_e2d4d651),
    .d(al_4caca369[0]),
    .o(al_186881f4));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_49199767 (
    .a(al_186881f4),
    .b(al_e31889d8[0]),
    .c(al_e31889d8[1]),
    .o(al_def29dc7));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_133614e6 (
    .a(al_def29dc7),
    .b(al_6db5b9d2),
    .c(al_e31889d8[2]),
    .d(al_e31889d8[3]),
    .e(al_e31889d8[4]),
    .o(al_322f98e5));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_389e140f (
    .a(al_def29dc7),
    .b(al_6db5b9d2),
    .c(al_e31889d8[2]),
    .d(al_e31889d8[3]),
    .o(al_45ef6b15));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_4e2adda6 (
    .a(al_186881f4),
    .b(al_6db5b9d2),
    .c(al_e31889d8[0]),
    .o(al_c3b5911e));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_b67e893 (
    .a(al_186881f4),
    .b(al_6db5b9d2),
    .c(al_e31889d8[0]),
    .d(al_e31889d8[1]),
    .o(al_e9d8781));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_e6c57e82 (
    .a(al_def29dc7),
    .b(al_6db5b9d2),
    .c(al_e31889d8[2]),
    .o(al_552a02c8));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_be3bdfea (
    .a(al_def29dc7),
    .b(al_6db5b9d2),
    .c(al_e31889d8[2]),
    .d(al_e31889d8[3]),
    .e(al_e31889d8[4]),
    .f(al_e31889d8[5]),
    .o(al_2684592f));
  AL_DFF_0 al_cc4859e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3b5911e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e31889d8[0]));
  AL_DFF_0 al_c92e567a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e9d8781),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e31889d8[1]));
  AL_DFF_0 al_905896d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_56ab2c31),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8349e0d1[2]));
  AL_DFF_0 al_18f667d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fdc5c136),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8349e0d1[3]));
  AL_DFF_0 al_51c621d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f838789f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8349e0d1[4]));
  AL_DFF_0 al_2e8aed30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_31c210),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8349e0d1[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_40b383f3 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_8349e0d1[0]),
    .e(al_8349e0d1[1]),
    .f(al_8349e0d1[2]),
    .o(al_e2323e1d));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_d7583022 (
    .a(al_e2323e1d),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_8349e0d1[3]),
    .f(al_8349e0d1[4]),
    .o(al_1b504c84));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_2f3afd0f (
    .a(al_1b504c84),
    .b(al_8349e0d1[5]),
    .c(al_5be1fa83),
    .d(al_b065182c[0]),
    .o(al_36b0c0a));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_6609f560 (
    .a(al_36b0c0a),
    .b(al_8349e0d1[0]),
    .c(al_8349e0d1[1]),
    .o(al_a201d3b2));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_a098a524 (
    .a(al_a201d3b2),
    .b(al_6db5b9d2),
    .c(al_8349e0d1[2]),
    .d(al_8349e0d1[3]),
    .e(al_8349e0d1[4]),
    .o(al_f838789f));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_d1a44480 (
    .a(al_a201d3b2),
    .b(al_6db5b9d2),
    .c(al_8349e0d1[2]),
    .d(al_8349e0d1[3]),
    .o(al_fdc5c136));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_a407bafd (
    .a(al_36b0c0a),
    .b(al_6db5b9d2),
    .c(al_8349e0d1[0]),
    .o(al_12797435));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_ebdc35b5 (
    .a(al_36b0c0a),
    .b(al_6db5b9d2),
    .c(al_8349e0d1[0]),
    .d(al_8349e0d1[1]),
    .o(al_eb32138));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_2d212cf1 (
    .a(al_a201d3b2),
    .b(al_6db5b9d2),
    .c(al_8349e0d1[2]),
    .o(al_56ab2c31));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_16f7d25d (
    .a(al_a201d3b2),
    .b(al_6db5b9d2),
    .c(al_8349e0d1[2]),
    .d(al_8349e0d1[3]),
    .e(al_8349e0d1[4]),
    .f(al_8349e0d1[5]),
    .o(al_31c210));
  AL_DFF_0 al_b73fd066 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_12797435),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8349e0d1[0]));
  AL_DFF_0 al_f442c9a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eb32138),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8349e0d1[1]));
  AL_DFF_0 al_80f6873e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_81f7233),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ef171e7[2]));
  AL_DFF_0 al_37137823 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_71703480),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ef171e7[3]));
  AL_DFF_0 al_879f4fb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d7bd990b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ef171e7[4]));
  AL_DFF_0 al_172756fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_739cb624),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ef171e7[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_8ff9a34 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_2ef171e7[0]),
    .e(al_2ef171e7[1]),
    .f(al_2ef171e7[2]),
    .o(al_73e64072));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_fec1a757 (
    .a(al_73e64072),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_2ef171e7[3]),
    .f(al_2ef171e7[4]),
    .o(al_84ac14c0));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_9882d9a0 (
    .a(al_84ac14c0),
    .b(al_2ef171e7[5]),
    .c(al_fd460907),
    .d(al_28515a17[0]),
    .o(al_eeb27c9c));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_e1a4ea35 (
    .a(al_eeb27c9c),
    .b(al_2ef171e7[0]),
    .c(al_2ef171e7[1]),
    .o(al_32cf3ccd));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_8bc932aa (
    .a(al_32cf3ccd),
    .b(al_6db5b9d2),
    .c(al_2ef171e7[2]),
    .d(al_2ef171e7[3]),
    .e(al_2ef171e7[4]),
    .o(al_d7bd990b));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_738b6e4f (
    .a(al_32cf3ccd),
    .b(al_6db5b9d2),
    .c(al_2ef171e7[2]),
    .d(al_2ef171e7[3]),
    .o(al_71703480));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_c83ab1a (
    .a(al_eeb27c9c),
    .b(al_6db5b9d2),
    .c(al_2ef171e7[0]),
    .o(al_9a4d5ae0));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_78c07ec5 (
    .a(al_eeb27c9c),
    .b(al_6db5b9d2),
    .c(al_2ef171e7[0]),
    .d(al_2ef171e7[1]),
    .o(al_6bb6f9ee));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_319633a5 (
    .a(al_32cf3ccd),
    .b(al_6db5b9d2),
    .c(al_2ef171e7[2]),
    .o(al_81f7233));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_a825863c (
    .a(al_32cf3ccd),
    .b(al_6db5b9d2),
    .c(al_2ef171e7[2]),
    .d(al_2ef171e7[3]),
    .e(al_2ef171e7[4]),
    .f(al_2ef171e7[5]),
    .o(al_739cb624));
  AL_DFF_0 al_abc4fc37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9a4d5ae0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ef171e7[0]));
  AL_DFF_0 al_df86823f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6bb6f9ee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ef171e7[1]));
  AL_DFF_0 al_3a2de498 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ea7f7c64),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_662b3089[2]));
  AL_DFF_0 al_deae4f28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80d96d10),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_662b3089[3]));
  AL_DFF_0 al_9850dc78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a98f5d5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_662b3089[4]));
  AL_DFF_0 al_b846e740 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_696ce813),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_662b3089[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_685605bb (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_662b3089[0]),
    .e(al_662b3089[1]),
    .f(al_662b3089[2]),
    .o(al_bd522ea7));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_97eecd68 (
    .a(al_bd522ea7),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_662b3089[3]),
    .f(al_662b3089[4]),
    .o(al_6aad2723));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_b4859e94 (
    .a(al_6aad2723),
    .b(al_662b3089[5]),
    .c(al_8815304a),
    .d(al_4caca369[0]),
    .o(al_422c6d68));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_eda0bd73 (
    .a(al_422c6d68),
    .b(al_662b3089[0]),
    .c(al_662b3089[1]),
    .o(al_aec0250a));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_5c4774cf (
    .a(al_aec0250a),
    .b(al_6db5b9d2),
    .c(al_662b3089[2]),
    .d(al_662b3089[3]),
    .e(al_662b3089[4]),
    .o(al_a98f5d5));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_4b12de46 (
    .a(al_aec0250a),
    .b(al_6db5b9d2),
    .c(al_662b3089[2]),
    .d(al_662b3089[3]),
    .o(al_80d96d10));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_29029fe9 (
    .a(al_422c6d68),
    .b(al_6db5b9d2),
    .c(al_662b3089[0]),
    .o(al_bcb724be));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_8f004d38 (
    .a(al_422c6d68),
    .b(al_6db5b9d2),
    .c(al_662b3089[0]),
    .d(al_662b3089[1]),
    .o(al_581cf91a));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_d03274e9 (
    .a(al_aec0250a),
    .b(al_6db5b9d2),
    .c(al_662b3089[2]),
    .o(al_ea7f7c64));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_9e9b175b (
    .a(al_aec0250a),
    .b(al_6db5b9d2),
    .c(al_662b3089[2]),
    .d(al_662b3089[3]),
    .e(al_662b3089[4]),
    .f(al_662b3089[5]),
    .o(al_696ce813));
  AL_DFF_0 al_9f8159bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bcb724be),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_662b3089[0]));
  AL_DFF_0 al_99faa371 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_581cf91a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_662b3089[1]));
  AL_DFF_0 al_19b0627e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2039287b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a30bd0f[2]));
  AL_DFF_0 al_c3123887 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_890d7ece),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a30bd0f[3]));
  AL_DFF_0 al_f0f0cae4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_290e28a2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a30bd0f[4]));
  AL_DFF_0 al_c0ac4587 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef0a54ec),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a30bd0f[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_2ffce6c (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_4a30bd0f[0]),
    .e(al_4a30bd0f[1]),
    .f(al_4a30bd0f[2]),
    .o(al_792502fb));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_455ad153 (
    .a(al_792502fb),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_4a30bd0f[3]),
    .f(al_4a30bd0f[4]),
    .o(al_fdf8d449));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_c8e305f9 (
    .a(al_fdf8d449),
    .b(al_4a30bd0f[5]),
    .c(al_2e8aa91),
    .d(al_4caca369[0]),
    .o(al_a540be99));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_26dea2fd (
    .a(al_a540be99),
    .b(al_4a30bd0f[0]),
    .c(al_4a30bd0f[1]),
    .d(al_4a30bd0f[2]),
    .e(al_4a30bd0f[3]),
    .f(al_4a30bd0f[4]),
    .o(al_34ca0b86));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_d9dbe655 (
    .a(al_a540be99),
    .b(al_4a30bd0f[0]),
    .c(al_4a30bd0f[1]),
    .d(al_4a30bd0f[2]),
    .e(al_4a30bd0f[3]),
    .f(al_4a30bd0f[4]),
    .o(al_90969885));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_99db7c2c (
    .a(al_90969885),
    .b(al_6db5b9d2),
    .o(al_290e28a2));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_2510cb6c (
    .a(al_a540be99),
    .b(al_6db5b9d2),
    .c(al_4a30bd0f[0]),
    .d(al_4a30bd0f[1]),
    .e(al_4a30bd0f[2]),
    .f(al_4a30bd0f[3]),
    .o(al_890d7ece));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_2be7cb8e (
    .a(al_a540be99),
    .b(al_6db5b9d2),
    .c(al_4a30bd0f[0]),
    .o(al_5fe1070b));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_2a2fcf8d (
    .a(al_a540be99),
    .b(al_6db5b9d2),
    .c(al_4a30bd0f[0]),
    .d(al_4a30bd0f[1]),
    .o(al_83fb54f8));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_c7ae2e6 (
    .a(al_a540be99),
    .b(al_6db5b9d2),
    .c(al_4a30bd0f[0]),
    .d(al_4a30bd0f[1]),
    .e(al_4a30bd0f[2]),
    .o(al_2039287b));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_195a37f9 (
    .a(al_34ca0b86),
    .b(al_6db5b9d2),
    .c(al_4a30bd0f[5]),
    .o(al_ef0a54ec));
  AL_DFF_0 al_a48b9ddf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5fe1070b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a30bd0f[0]));
  AL_DFF_0 al_6f5932cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_83fb54f8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a30bd0f[1]));
  AL_DFF_0 al_fe6e92b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d44a1539),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2119f32d[2]));
  AL_DFF_0 al_e1ac7b7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5e34a0d9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2119f32d[3]));
  AL_DFF_0 al_89f06a5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_187efcc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2119f32d[4]));
  AL_DFF_0 al_ea8dfa0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_691042b7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2119f32d[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_e3ee5571 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_2119f32d[0]),
    .e(al_2119f32d[1]),
    .f(al_2119f32d[2]),
    .o(al_eefb494d));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_3c0489ae (
    .a(al_eefb494d),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_2119f32d[3]),
    .f(al_2119f32d[4]),
    .o(al_733e11d7));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_70a828bb (
    .a(al_733e11d7),
    .b(al_2119f32d[5]),
    .c(al_ce1c71c5),
    .d(al_b065182c[0]),
    .o(al_eb9d8684));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_daf432f9 (
    .a(al_eb9d8684),
    .b(al_2119f32d[0]),
    .c(al_2119f32d[1]),
    .o(al_9e7f07bf));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_cb698127 (
    .a(al_9e7f07bf),
    .b(al_6db5b9d2),
    .c(al_2119f32d[2]),
    .d(al_2119f32d[3]),
    .e(al_2119f32d[4]),
    .o(al_187efcc));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_38b553d (
    .a(al_9e7f07bf),
    .b(al_6db5b9d2),
    .c(al_2119f32d[2]),
    .d(al_2119f32d[3]),
    .o(al_5e34a0d9));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_49c817f1 (
    .a(al_eb9d8684),
    .b(al_6db5b9d2),
    .c(al_2119f32d[0]),
    .o(al_70337de1));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_be452956 (
    .a(al_eb9d8684),
    .b(al_6db5b9d2),
    .c(al_2119f32d[0]),
    .d(al_2119f32d[1]),
    .o(al_da48a4d6));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_9f757af4 (
    .a(al_9e7f07bf),
    .b(al_6db5b9d2),
    .c(al_2119f32d[2]),
    .o(al_d44a1539));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_42e220a0 (
    .a(al_9e7f07bf),
    .b(al_6db5b9d2),
    .c(al_2119f32d[2]),
    .d(al_2119f32d[3]),
    .e(al_2119f32d[4]),
    .f(al_2119f32d[5]),
    .o(al_691042b7));
  AL_DFF_0 al_df0f883b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_70337de1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2119f32d[0]));
  AL_DFF_0 al_f88f856e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_da48a4d6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2119f32d[1]));
  AL_DFF_0 al_54c5c843 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f6e3dfbd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9591ec3[2]));
  AL_DFF_0 al_2efebb35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_810f7f51),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9591ec3[3]));
  AL_DFF_0 al_91bce73d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3077309),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9591ec3[4]));
  AL_DFF_0 al_efe53875 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ff2cde7a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9591ec3[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_c28acd85 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_d9591ec3[0]),
    .e(al_d9591ec3[1]),
    .f(al_d9591ec3[2]),
    .o(al_c0cdd2f2));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_a963936f (
    .a(al_c0cdd2f2),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_d9591ec3[3]),
    .f(al_d9591ec3[4]),
    .o(al_3ed1abca));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_71c7056a (
    .a(al_3ed1abca),
    .b(al_d9591ec3[5]),
    .c(al_9929d21),
    .d(al_28515a17[0]),
    .o(al_31adef42));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_3de5873a (
    .a(al_31adef42),
    .b(al_d9591ec3[0]),
    .c(al_d9591ec3[1]),
    .o(al_223e27a1));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_b1d2433e (
    .a(al_223e27a1),
    .b(al_6db5b9d2),
    .c(al_d9591ec3[2]),
    .d(al_d9591ec3[3]),
    .e(al_d9591ec3[4]),
    .o(al_c3077309));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_870b7fca (
    .a(al_223e27a1),
    .b(al_6db5b9d2),
    .c(al_d9591ec3[2]),
    .d(al_d9591ec3[3]),
    .o(al_810f7f51));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_f1add8b7 (
    .a(al_31adef42),
    .b(al_6db5b9d2),
    .c(al_d9591ec3[0]),
    .o(al_6224ca70));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_c8a0e4f4 (
    .a(al_31adef42),
    .b(al_6db5b9d2),
    .c(al_d9591ec3[0]),
    .d(al_d9591ec3[1]),
    .o(al_77706154));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_a83d724c (
    .a(al_223e27a1),
    .b(al_6db5b9d2),
    .c(al_d9591ec3[2]),
    .o(al_f6e3dfbd));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_8d6e2cd4 (
    .a(al_223e27a1),
    .b(al_6db5b9d2),
    .c(al_d9591ec3[2]),
    .d(al_d9591ec3[3]),
    .e(al_d9591ec3[4]),
    .f(al_d9591ec3[5]),
    .o(al_ff2cde7a));
  AL_DFF_0 al_7906588d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6224ca70),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9591ec3[0]));
  AL_DFF_0 al_a4fa4ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_77706154),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9591ec3[1]));
  AL_DFF_0 al_c444aad8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d6502391),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_ee7571b0));
  AL_DFF_0 al_a39fa0d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_89b57934),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_b0c5cb0b));
  AL_DFF_0 al_760e0b1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ce868614),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_b09b809));
  AL_DFF_0 al_a9404307 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6a0200a0),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_ba71435f));
  AL_DFF_0 al_a5629b51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d93c50d7),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_b40c9ab5));
  AL_DFF_0 al_6f4b350d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2ebef479),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_fbbf0c04));
  AL_DFF_0 al_95e7c800 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4cb605a3),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_335c3c71));
  AL_DFF_0 al_e16409c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3f7b50be),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_be14e3f3));
  AL_DFF_0 al_170e40f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4531bc64),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_31cf7bc9));
  AL_DFF_0 al_7b7b0809 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9b495b9),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_8e660235));
  AL_DFF_0 al_5f86cee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_472a7b46),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_e6d4af1));
  AL_DFF_0 al_6c878b42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bf50c51c),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_1759a3a0));
  AL_DFF_0 al_e015aff6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a07095e8),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_30c9bd77));
  AL_DFF_0 al_3e003084 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3b280eeb),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_6f07b96e));
  AL_DFF_0 al_5e56e66e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b4d25a49),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_4ab9f9ad));
  AL_DFF_0 al_782d8468 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_92250858),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7c6973e));
  AL_DFF_0 al_95b7bc29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3f68feff),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_1f596d24));
  AL_DFF_0 al_281e6513 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a7a585be),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_dc57999f));
  AL_DFF_0 al_f64f683c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef6d9f73),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_f9e69b00));
  AL_DFF_0 al_f7cba562 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b285e414),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_3a2d553d));
  AL_DFF_0 al_d19f5ce0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4783da3f),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_a88d3bd8));
  AL_DFF_0 al_c7b941dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f45ad02a),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_722c0dcd));
  AL_DFF_0 al_50e02094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_130738c8),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_4e018b61));
  AL_DFF_0 al_30c9b643 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_14656fdb),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_1f414bbe));
  AL_DFF_0 al_bc3cc471 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f9fd3044),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_eadb4e14));
  AL_DFF_0 al_8a569ada (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1abf75fc),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_a771a309));
  AL_DFF_0 al_427c75bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ee3904b1),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_20f5f77c));
  AL_DFF_0 al_bd771ac1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_96b7453),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_d88aee38));
  AL_DFF_0 al_bee17a08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3858b210),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_f9c30b23));
  AL_DFF_0 al_4e297471 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55b9d73d),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_d2a2bf32));
  AL_DFF_0 al_df90a296 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6f9c4eba),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_c41fccfb));
  AL_DFF_0 al_93acd318 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_664e4e8f),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_91458dff));
  AL_DFF_0 al_b34456e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_852588b2),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_ade031de));
  AL_DFF_0 al_e3e4d20d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_14200974),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_830e948));
  AL_DFF_0 al_3beebd0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f3b50940),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_d0276689));
  AL_DFF_0 al_e4c18951 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_da329b96),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_8e003744));
  AL_DFF_0 al_e68d586b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ca5b293f),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_8d08d03c));
  AL_DFF_0 al_15504ae9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b57594f0),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_e470f61d));
  AL_DFF_0 al_aee65fcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_15554a76),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_93161d1e));
  AL_DFF_0 al_3b755c40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e3bba389),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_77d022d8));
  AL_DFF_0 al_1c85fb23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cda79e31),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_c732c324));
  AL_DFF_0 al_2cbfea5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7aee3607),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_fbdc3092));
  AL_DFF_0 al_ad4d9741 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9a683f3),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_142dd1c8));
  AL_DFF_0 al_9b6172b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_80baf9fa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d102248[2]));
  AL_DFF_0 al_45536fc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c9b8e286),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d102248[3]));
  AL_DFF_0 al_6b5dd4e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7038cb56),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d102248[4]));
  AL_DFF_0 al_ee43b11f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_309702b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d102248[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_bf9cab70 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_1d102248[0]),
    .e(al_1d102248[1]),
    .f(al_1d102248[2]),
    .o(al_61b9dbed));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_9d947b0 (
    .a(al_61b9dbed),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_1d102248[3]),
    .f(al_1d102248[4]),
    .o(al_27d43db3));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_4f3bdade (
    .a(al_27d43db3),
    .b(al_1d102248[5]),
    .c(al_23ce284b),
    .d(al_4caca369[0]),
    .o(al_401f1215));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_cca6f5b2 (
    .a(al_401f1215),
    .b(al_1d102248[0]),
    .c(al_1d102248[1]),
    .d(al_1d102248[2]),
    .e(al_1d102248[3]),
    .f(al_1d102248[4]),
    .o(al_5d0bc72b));
  AL_MAP_LUT6 #(
    .EQN("~(F@(E*D*C*B*~A))"),
    .INIT(64'h40000000bfffffff))
    al_75dbe573 (
    .a(al_401f1215),
    .b(al_1d102248[0]),
    .c(al_1d102248[1]),
    .d(al_1d102248[2]),
    .e(al_1d102248[3]),
    .f(al_1d102248[4]),
    .o(al_ad7bbe14));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_d2d7d86e (
    .a(al_ad7bbe14),
    .b(al_6db5b9d2),
    .o(al_7038cb56));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_e3b9ce10 (
    .a(al_401f1215),
    .b(al_6db5b9d2),
    .c(al_1d102248[0]),
    .d(al_1d102248[1]),
    .e(al_1d102248[2]),
    .f(al_1d102248[3]),
    .o(al_c9b8e286));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_59306353 (
    .a(al_401f1215),
    .b(al_6db5b9d2),
    .c(al_1d102248[0]),
    .o(al_a0a71833));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_1de0a75d (
    .a(al_401f1215),
    .b(al_6db5b9d2),
    .c(al_1d102248[0]),
    .d(al_1d102248[1]),
    .o(al_9cc84a67));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_78f62c04 (
    .a(al_401f1215),
    .b(al_6db5b9d2),
    .c(al_1d102248[0]),
    .d(al_1d102248[1]),
    .e(al_1d102248[2]),
    .o(al_80baf9fa));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_a3ee0d4b (
    .a(al_5d0bc72b),
    .b(al_6db5b9d2),
    .c(al_1d102248[5]),
    .o(al_309702b));
  AL_DFF_0 al_1c88d501 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a0a71833),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d102248[0]));
  AL_DFF_0 al_1ff23661 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9cc84a67),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d102248[1]));
  AL_DFF_0 al_aab47c15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dac9476c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f78383db[2]));
  AL_DFF_0 al_b9431ed7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2f7efa54),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f78383db[3]));
  AL_DFF_0 al_ae42ff20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_85e91cf0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f78383db[4]));
  AL_DFF_0 al_6bcf6ef9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_527ad770),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f78383db[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_c791d3c (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_f78383db[0]),
    .e(al_f78383db[1]),
    .f(al_f78383db[2]),
    .o(al_e4e2df3a));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_6745ef4d (
    .a(al_e4e2df3a),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_f78383db[3]),
    .f(al_f78383db[4]),
    .o(al_e1d70a3d));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_2879b47d (
    .a(al_e1d70a3d),
    .b(al_f78383db[5]),
    .c(al_4aba11ac),
    .d(al_b065182c[0]),
    .o(al_50c08ac));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_36519d72 (
    .a(al_50c08ac),
    .b(al_f78383db[0]),
    .c(al_f78383db[1]),
    .o(al_163e3e0c));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_bd1a2ae3 (
    .a(al_163e3e0c),
    .b(al_6db5b9d2),
    .c(al_f78383db[2]),
    .d(al_f78383db[3]),
    .e(al_f78383db[4]),
    .o(al_85e91cf0));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_36409aa8 (
    .a(al_163e3e0c),
    .b(al_6db5b9d2),
    .c(al_f78383db[2]),
    .d(al_f78383db[3]),
    .o(al_2f7efa54));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_aeecca77 (
    .a(al_50c08ac),
    .b(al_6db5b9d2),
    .c(al_f78383db[0]),
    .o(al_bbb63b9));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_64a0cd0d (
    .a(al_50c08ac),
    .b(al_6db5b9d2),
    .c(al_f78383db[0]),
    .d(al_f78383db[1]),
    .o(al_e4a5394c));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_4d861645 (
    .a(al_163e3e0c),
    .b(al_6db5b9d2),
    .c(al_f78383db[2]),
    .o(al_dac9476c));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_70b36ee9 (
    .a(al_163e3e0c),
    .b(al_6db5b9d2),
    .c(al_f78383db[2]),
    .d(al_f78383db[3]),
    .e(al_f78383db[4]),
    .f(al_f78383db[5]),
    .o(al_527ad770));
  AL_DFF_0 al_c7734a48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bbb63b9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f78383db[0]));
  AL_DFF_0 al_9cc24bbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e4a5394c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f78383db[1]));
  AL_DFF_0 al_64b33dcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1556ef5b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9be1f39[2]));
  AL_DFF_0 al_2876000e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e0f76854),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9be1f39[3]));
  AL_DFF_0 al_b693d126 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bbd8d9ee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9be1f39[4]));
  AL_DFF_0 al_c76134fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9f44cd3f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9be1f39[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_f5395dd4 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_d9be1f39[0]),
    .e(al_d9be1f39[1]),
    .f(al_d9be1f39[2]),
    .o(al_bd9db94a));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_a22dfbf5 (
    .a(al_bd9db94a),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_d9be1f39[3]),
    .f(al_d9be1f39[4]),
    .o(al_898acbc2));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_c0418d9b (
    .a(al_898acbc2),
    .b(al_d9be1f39[5]),
    .c(al_20c1f74d),
    .d(al_28515a17[0]),
    .o(al_81777b16));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_d6c4ca4e (
    .a(al_81777b16),
    .b(al_d9be1f39[0]),
    .c(al_d9be1f39[1]),
    .d(al_d9be1f39[2]),
    .e(al_d9be1f39[3]),
    .f(al_d9be1f39[4]),
    .o(al_f996058d));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_54f9f644 (
    .a(al_81777b16),
    .b(al_d9be1f39[0]),
    .c(al_d9be1f39[1]),
    .d(al_d9be1f39[2]),
    .e(al_d9be1f39[3]),
    .f(al_d9be1f39[4]),
    .o(al_7fda6214));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_e486d4d6 (
    .a(al_7fda6214),
    .b(al_6db5b9d2),
    .o(al_bbd8d9ee));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_60a8ea63 (
    .a(al_81777b16),
    .b(al_6db5b9d2),
    .c(al_d9be1f39[0]),
    .d(al_d9be1f39[1]),
    .e(al_d9be1f39[2]),
    .f(al_d9be1f39[3]),
    .o(al_e0f76854));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_bb8cbae (
    .a(al_81777b16),
    .b(al_6db5b9d2),
    .c(al_d9be1f39[0]),
    .o(al_d524c6a5));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_5fd8ade1 (
    .a(al_81777b16),
    .b(al_6db5b9d2),
    .c(al_d9be1f39[0]),
    .d(al_d9be1f39[1]),
    .o(al_a6968310));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_ffe5a29d (
    .a(al_81777b16),
    .b(al_6db5b9d2),
    .c(al_d9be1f39[0]),
    .d(al_d9be1f39[1]),
    .e(al_d9be1f39[2]),
    .o(al_1556ef5b));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_22897e07 (
    .a(al_f996058d),
    .b(al_6db5b9d2),
    .c(al_d9be1f39[5]),
    .o(al_9f44cd3f));
  AL_DFF_0 al_5e7fa70e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d524c6a5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9be1f39[0]));
  AL_DFF_0 al_62aff4fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a6968310),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d9be1f39[1]));
  AL_DFF_0 al_7f96e615 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7bd1a9d6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e255230[2]));
  AL_DFF_0 al_dc5b2da8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_31b57a77),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e255230[3]));
  AL_DFF_0 al_e8545e9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c3f3285c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e255230[4]));
  AL_DFF_0 al_a249300c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7d2b45a1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e255230[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_85dbad5a (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_1e255230[0]),
    .e(al_1e255230[1]),
    .f(al_1e255230[2]),
    .o(al_2fdd1128));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_84c1accf (
    .a(al_2fdd1128),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_1e255230[3]),
    .f(al_1e255230[4]),
    .o(al_6d6f3341));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_974e8a83 (
    .a(al_6d6f3341),
    .b(al_1e255230[5]),
    .c(al_8fa72152),
    .d(al_4caca369[0]),
    .o(al_fbacc3a8));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_2d4a0377 (
    .a(al_fbacc3a8),
    .b(al_1e255230[0]),
    .c(al_1e255230[1]),
    .o(al_b9053852));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_6976f9ed (
    .a(al_b9053852),
    .b(al_6db5b9d2),
    .c(al_1e255230[2]),
    .d(al_1e255230[3]),
    .e(al_1e255230[4]),
    .o(al_c3f3285c));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_715c169c (
    .a(al_b9053852),
    .b(al_6db5b9d2),
    .c(al_1e255230[2]),
    .d(al_1e255230[3]),
    .o(al_31b57a77));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_fbcde7f8 (
    .a(al_fbacc3a8),
    .b(al_6db5b9d2),
    .c(al_1e255230[0]),
    .o(al_f1d76027));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_f253ef05 (
    .a(al_fbacc3a8),
    .b(al_6db5b9d2),
    .c(al_1e255230[0]),
    .d(al_1e255230[1]),
    .o(al_cdb85e5d));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_1d3e5861 (
    .a(al_b9053852),
    .b(al_6db5b9d2),
    .c(al_1e255230[2]),
    .o(al_7bd1a9d6));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_d5fd70e5 (
    .a(al_b9053852),
    .b(al_6db5b9d2),
    .c(al_1e255230[2]),
    .d(al_1e255230[3]),
    .e(al_1e255230[4]),
    .f(al_1e255230[5]),
    .o(al_7d2b45a1));
  AL_DFF_0 al_f898b651 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f1d76027),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e255230[0]));
  AL_DFF_0 al_c850618d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cdb85e5d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1e255230[1]));
  AL_DFF_0 al_b14f25e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_312f6ab1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d61bccef[2]));
  AL_DFF_0 al_31447466 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7b6b3d00),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d61bccef[3]));
  AL_DFF_0 al_3efdc824 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b349d1f9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d61bccef[4]));
  AL_DFF_0 al_579b0961 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_241ce585),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d61bccef[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_ad4b4c60 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_d61bccef[0]),
    .e(al_d61bccef[1]),
    .f(al_d61bccef[2]),
    .o(al_3f1b9f0e));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_27b4e877 (
    .a(al_3f1b9f0e),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_d61bccef[3]),
    .f(al_d61bccef[4]),
    .o(al_316d230a));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_3287b368 (
    .a(al_316d230a),
    .b(al_d61bccef[5]),
    .c(al_ea6ecc89),
    .d(al_b065182c[0]),
    .o(al_8b91849a));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_dfbe594f (
    .a(al_8b91849a),
    .b(al_d61bccef[0]),
    .c(al_d61bccef[1]),
    .o(al_e220508d));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_2846ef61 (
    .a(al_e220508d),
    .b(al_6db5b9d2),
    .c(al_d61bccef[2]),
    .d(al_d61bccef[3]),
    .e(al_d61bccef[4]),
    .o(al_b349d1f9));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_fb8f3ce8 (
    .a(al_e220508d),
    .b(al_6db5b9d2),
    .c(al_d61bccef[2]),
    .d(al_d61bccef[3]),
    .o(al_7b6b3d00));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_b4c0c46e (
    .a(al_8b91849a),
    .b(al_6db5b9d2),
    .c(al_d61bccef[0]),
    .o(al_5fc98ca9));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_692528b2 (
    .a(al_8b91849a),
    .b(al_6db5b9d2),
    .c(al_d61bccef[0]),
    .d(al_d61bccef[1]),
    .o(al_e42e193d));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_5d2452d4 (
    .a(al_e220508d),
    .b(al_6db5b9d2),
    .c(al_d61bccef[2]),
    .o(al_312f6ab1));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_ee84be3b (
    .a(al_e220508d),
    .b(al_6db5b9d2),
    .c(al_d61bccef[2]),
    .d(al_d61bccef[3]),
    .e(al_d61bccef[4]),
    .f(al_d61bccef[5]),
    .o(al_241ce585));
  AL_DFF_0 al_c74a63d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5fc98ca9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d61bccef[0]));
  AL_DFF_0 al_c7f0eab0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e42e193d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d61bccef[1]));
  AL_DFF_0 al_3d91002a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c4ec8088),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46e8788c[2]));
  AL_DFF_0 al_1a7f59cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7a2b0bb8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46e8788c[3]));
  AL_DFF_0 al_83731a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ebe8b3b7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46e8788c[4]));
  AL_DFF_0 al_a4cfd6e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_920bfd47),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46e8788c[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_4745bcc0 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_46e8788c[0]),
    .e(al_46e8788c[1]),
    .f(al_46e8788c[2]),
    .o(al_54647363));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_9580380a (
    .a(al_54647363),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_46e8788c[3]),
    .f(al_46e8788c[4]),
    .o(al_e75d67c1));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_e4c73127 (
    .a(al_e75d67c1),
    .b(al_46e8788c[5]),
    .c(al_10f5be33),
    .d(al_28515a17[0]),
    .o(al_fbdfd137));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_e85045f1 (
    .a(al_fbdfd137),
    .b(al_46e8788c[0]),
    .c(al_46e8788c[1]),
    .o(al_b10901c4));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_572fc0e7 (
    .a(al_b10901c4),
    .b(al_6db5b9d2),
    .c(al_46e8788c[2]),
    .d(al_46e8788c[3]),
    .e(al_46e8788c[4]),
    .o(al_ebe8b3b7));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_2f95c82 (
    .a(al_b10901c4),
    .b(al_6db5b9d2),
    .c(al_46e8788c[2]),
    .d(al_46e8788c[3]),
    .o(al_7a2b0bb8));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_fae8f8a7 (
    .a(al_fbdfd137),
    .b(al_6db5b9d2),
    .c(al_46e8788c[0]),
    .o(al_ba559767));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_53f16d2a (
    .a(al_fbdfd137),
    .b(al_6db5b9d2),
    .c(al_46e8788c[0]),
    .d(al_46e8788c[1]),
    .o(al_189beaf8));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_3d221f61 (
    .a(al_b10901c4),
    .b(al_6db5b9d2),
    .c(al_46e8788c[2]),
    .o(al_c4ec8088));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_57b8b4b1 (
    .a(al_b10901c4),
    .b(al_6db5b9d2),
    .c(al_46e8788c[2]),
    .d(al_46e8788c[3]),
    .e(al_46e8788c[4]),
    .f(al_46e8788c[5]),
    .o(al_920bfd47));
  AL_DFF_0 al_af172ac8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ba559767),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46e8788c[0]));
  AL_DFF_0 al_c9f6b6b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_189beaf8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46e8788c[1]));
  AL_DFF_0 al_1bda7a8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d2207ab),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56e72bf4[2]));
  AL_DFF_0 al_9a7275f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b7580b14),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56e72bf4[3]));
  AL_DFF_0 al_81f63cb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_84c4e89e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56e72bf4[4]));
  AL_DFF_0 al_5d91a37c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4e77858f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56e72bf4[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_2e8011ee (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_56e72bf4[0]),
    .e(al_56e72bf4[1]),
    .f(al_56e72bf4[2]),
    .o(al_b627b129));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_433f4bf7 (
    .a(al_b627b129),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_56e72bf4[3]),
    .f(al_56e72bf4[4]),
    .o(al_ec10e78f));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_55b2af36 (
    .a(al_ec10e78f),
    .b(al_56e72bf4[5]),
    .c(al_d90f1fe1),
    .d(al_4caca369[0]),
    .o(al_c4cdc14c));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_a953c30f (
    .a(al_c4cdc14c),
    .b(al_56e72bf4[0]),
    .c(al_56e72bf4[1]),
    .o(al_c88a646f));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_7576edcc (
    .a(al_c88a646f),
    .b(al_6db5b9d2),
    .c(al_56e72bf4[2]),
    .d(al_56e72bf4[3]),
    .e(al_56e72bf4[4]),
    .o(al_84c4e89e));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_5867a9c7 (
    .a(al_c88a646f),
    .b(al_6db5b9d2),
    .c(al_56e72bf4[2]),
    .d(al_56e72bf4[3]),
    .o(al_b7580b14));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_3552c11c (
    .a(al_c4cdc14c),
    .b(al_6db5b9d2),
    .c(al_56e72bf4[0]),
    .o(al_d0e0cc74));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_f4272708 (
    .a(al_c4cdc14c),
    .b(al_6db5b9d2),
    .c(al_56e72bf4[0]),
    .d(al_56e72bf4[1]),
    .o(al_7077034d));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_a612a053 (
    .a(al_c88a646f),
    .b(al_6db5b9d2),
    .c(al_56e72bf4[2]),
    .o(al_4d2207ab));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_21596d1c (
    .a(al_c88a646f),
    .b(al_6db5b9d2),
    .c(al_56e72bf4[2]),
    .d(al_56e72bf4[3]),
    .e(al_56e72bf4[4]),
    .f(al_56e72bf4[5]),
    .o(al_4e77858f));
  AL_DFF_0 al_685993ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d0e0cc74),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56e72bf4[0]));
  AL_DFF_0 al_63199ca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7077034d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56e72bf4[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_52806057 (
    .a(al_6db5b9d2),
    .b(al_23ce284b),
    .c(al_6bddd01a),
    .o(al_748cb5ab));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_33b6f11f (
    .a(al_6db5b9d2),
    .b(al_9929d21),
    .c(al_83ebd977),
    .o(al_cc0caf5a));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_f7a0d861 (
    .a(al_6db5b9d2),
    .b(al_ce1c71c5),
    .c(al_c3e70575),
    .o(al_3f8224e9));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_d2928af2 (
    .a(al_6db5b9d2),
    .b(al_8815304a),
    .c(al_4864d933),
    .o(al_2534fd55));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_423d5a8b (
    .a(al_6db5b9d2),
    .b(al_fd460907),
    .c(al_4708b339),
    .o(al_de545759));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_2e4bf6d6 (
    .a(al_6db5b9d2),
    .b(al_5be1fa83),
    .c(al_2efa36ca),
    .o(al_aa84749f));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_4eec7c53 (
    .a(al_6db5b9d2),
    .b(al_e2d4d651),
    .c(al_5e6f3859),
    .o(al_1df0d799));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_82390141 (
    .a(al_6db5b9d2),
    .b(al_770f9dd1),
    .c(al_35f768f4),
    .o(al_421f3e11));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_a76785f5 (
    .a(al_6db5b9d2),
    .b(al_6e370c03),
    .c(al_ee615f87),
    .o(al_f06f70db));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_82cc98d (
    .a(al_6db5b9d2),
    .b(al_25e4ab96),
    .c(al_cc2e5bcc),
    .o(al_78d64c6e));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_423bc475 (
    .a(al_6db5b9d2),
    .b(al_7bafa36d),
    .c(al_31be1d74),
    .o(al_9898f5d2));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_df4fce96 (
    .a(al_6db5b9d2),
    .b(al_8b05cae6),
    .c(al_b56307ec),
    .o(al_3128e6f));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_a9f442ac (
    .a(al_6db5b9d2),
    .b(al_8dc56974),
    .c(al_7cd149c6),
    .o(al_a75ec498));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_b75bddf8 (
    .a(al_6db5b9d2),
    .b(al_1919cac5),
    .c(al_28d8d34d),
    .o(al_3c9faf77));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_1231f837 (
    .a(al_6db5b9d2),
    .b(al_521fd670),
    .c(al_a9490be8),
    .o(al_ce0ffb93));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_6f9bb246 (
    .a(al_6db5b9d2),
    .b(al_a48594d3),
    .c(al_9dcab982),
    .o(al_c2d49ea8));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_1b5698a1 (
    .a(al_6db5b9d2),
    .b(al_d27a1279),
    .c(al_2bb74c3d),
    .o(al_46e8cf64));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_780a17f0 (
    .a(al_6db5b9d2),
    .b(al_2fc8b96e),
    .c(al_80360204),
    .o(al_bfe09e38));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_2125f462 (
    .a(al_6db5b9d2),
    .b(al_8d8df5a3),
    .c(al_6dc98a03),
    .o(al_785b323e));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_eba5a7a6 (
    .a(al_6db5b9d2),
    .b(al_7bbb36d3),
    .c(al_df7aa915),
    .o(al_63db5a9c));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_77af6f98 (
    .a(al_6db5b9d2),
    .b(al_6db10ea9),
    .c(al_796e34c4),
    .o(al_98025056));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_16a029f (
    .a(al_6db5b9d2),
    .b(al_e2f3bed2),
    .c(al_fef4ecdb),
    .o(al_eaf1b77d));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_1138fda1 (
    .a(al_6db5b9d2),
    .b(al_24944e5c),
    .c(al_b8da0e9e),
    .o(al_64ae12a2));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_8ea744e5 (
    .a(al_6db5b9d2),
    .b(al_d4c409ba),
    .c(al_c81182c),
    .o(al_41c60d64));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_d05ff26 (
    .a(al_6db5b9d2),
    .b(al_4f9aa153),
    .c(al_ab1b2b16),
    .o(al_74787620));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_a8b807c0 (
    .a(al_6db5b9d2),
    .b(al_c9d182cf),
    .c(al_64f79045),
    .o(al_ef3dcd46));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_da43e26 (
    .a(al_6db5b9d2),
    .b(al_72ab91cb),
    .c(al_d9d76d0a),
    .o(al_956bd9e3));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_8091f81e (
    .a(al_6db5b9d2),
    .b(al_df90085e),
    .c(al_3da9562a),
    .o(al_82ccfd38));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_fb7e724e (
    .a(al_6db5b9d2),
    .b(al_17b42586),
    .c(al_21d51e65),
    .o(al_a9ba8e79));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_93a7ae20 (
    .a(al_6db5b9d2),
    .b(al_535f72cd),
    .c(al_9f6750b6),
    .o(al_17c12787));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_29112ccf (
    .a(al_6db5b9d2),
    .b(al_843f6bac),
    .c(al_82133c54),
    .o(al_5d326e5d));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_d72bdbc (
    .a(al_6db5b9d2),
    .b(al_87f40037),
    .c(al_106fddab),
    .o(al_b6bc6cf7));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_fc002748 (
    .a(al_6db5b9d2),
    .b(al_815c8034),
    .c(al_b8cc00cf),
    .o(al_caca8068));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_a3e62d52 (
    .a(al_6db5b9d2),
    .b(al_d90f1fe1),
    .c(al_12b38499),
    .o(al_ab39876a));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_fc2b4e70 (
    .a(al_6db5b9d2),
    .b(al_10f5be33),
    .c(al_3d66f550),
    .o(al_44b75b16));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_5c681817 (
    .a(al_6db5b9d2),
    .b(al_ea6ecc89),
    .c(al_ad58fbc9),
    .o(al_4359f728));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_53fe28ed (
    .a(al_6db5b9d2),
    .b(al_8fa72152),
    .c(al_ac593c94),
    .o(al_320b8e92));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_ac1305b7 (
    .a(al_6db5b9d2),
    .b(al_20c1f74d),
    .c(al_f7c9608b),
    .o(al_16e3e4ef));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_d0b30738 (
    .a(al_6db5b9d2),
    .b(al_4aba11ac),
    .c(al_c85cbcb),
    .o(al_9cb4bf74));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_5f702dad (
    .a(al_6db5b9d2),
    .b(al_2e8aa91),
    .c(al_71cac35e),
    .o(al_df8baf16));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_b245f1e8 (
    .a(al_6db5b9d2),
    .b(al_6e50ac65),
    .c(al_e6ea44e6),
    .o(al_881110e));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_ab30bdf3 (
    .a(al_6db5b9d2),
    .b(al_e2476620),
    .c(al_9b5a4dbd),
    .o(al_997d115c));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_7313b924 (
    .a(al_6db5b9d2),
    .b(al_9a6187ef),
    .c(al_4b4a698a),
    .o(al_b9ce4338));
  AL_DFF_0 al_77262bd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b9ce4338),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26a2c365));
  AL_DFF_0 al_e38c5dc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_997d115c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_55882f9d));
  AL_DFF_0 al_6b2d2112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_881110e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_267f05f8));
  AL_DFF_0 al_e7ff695a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_df8baf16),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c600a777));
  AL_DFF_0 al_c20a476c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9cb4bf74),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_435ecf83));
  AL_DFF_0 al_ded4ba74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_16e3e4ef),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c802abc3));
  AL_DFF_0 al_64be7edd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_320b8e92),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6615be3));
  AL_DFF_0 al_c85dd0f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4359f728),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53c183a7));
  AL_DFF_0 al_b6718f76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44b75b16),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b7e1c0f));
  AL_DFF_0 al_ff8378ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ab39876a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_228163ab));
  AL_DFF_0 al_137dd3c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_caca8068),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33cf56b3));
  AL_DFF_0 al_5bfd987f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b6bc6cf7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_39705b9f));
  AL_DFF_0 al_cc3e5f23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5d326e5d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_860bc871));
  AL_DFF_0 al_fb311279 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_17c12787),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eda53b41));
  AL_DFF_0 al_9f3b7655 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a9ba8e79),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8695553e));
  AL_DFF_0 al_b60a39a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_82ccfd38),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_646f260c));
  AL_DFF_0 al_11664bdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_956bd9e3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c63960b));
  AL_DFF_0 al_fa9bc53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ef3dcd46),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cea991a));
  AL_DFF_0 al_243fce59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_74787620),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fdd1bba3));
  AL_DFF_0 al_7f21fdc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41c60d64),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7ceaf80e));
  AL_DFF_0 al_a082bff3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_64ae12a2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_314e2528));
  AL_DFF_0 al_db0713ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_eaf1b77d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74f1ae6b));
  AL_DFF_0 al_4e7d1010 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_98025056),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49840bbd));
  AL_DFF_0 al_1020f42c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_63db5a9c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fa62f20b));
  AL_DFF_0 al_7da8af29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_785b323e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7da0d957));
  AL_DFF_0 al_d219c7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bfe09e38),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53b6ba74));
  AL_DFF_0 al_6cda4de0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46e8cf64),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46888ef2));
  AL_DFF_0 al_ea6c564b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c2d49ea8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c43abb));
  AL_DFF_0 al_994a8285 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ce0ffb93),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89f795c9));
  AL_DFF_0 al_4caf0f5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3c9faf77),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_652cea26));
  AL_DFF_0 al_43f5e1d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a75ec498),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f52bc7e));
  AL_DFF_0 al_fb5c7256 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3128e6f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14f4e684));
  AL_DFF_0 al_f4a919f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9898f5d2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1bbf8570));
  AL_DFF_0 al_298fe739 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_78d64c6e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59fdd957));
  AL_DFF_0 al_f6d07b3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f06f70db),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4e23dc54));
  AL_DFF_0 al_703b5fd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_421f3e11),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d79d15f2));
  AL_DFF_0 al_febceaed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1df0d799),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e956701b));
  AL_DFF_0 al_ac30aa85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aa84749f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3ec6ca0b));
  AL_DFF_0 al_ab07e17d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_de545759),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_38793d0));
  AL_DFF_0 al_48ffe3ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2534fd55),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3ea78ea2));
  AL_DFF_0 al_b4014f14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3f8224e9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c678f752));
  AL_DFF_0 al_8b0497ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cc0caf5a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5f1c8d24));
  AL_DFF_0 al_790053cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_748cb5ab),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ef6225f5));
  AL_DFF_0 al_b8f00388 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e49c184e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_620ff4d8[2]));
  AL_DFF_0 al_bea1456b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c958e833),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_620ff4d8[3]));
  AL_DFF_0 al_1c8c540a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3e72c22b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_620ff4d8[4]));
  AL_DFF_0 al_2736c4f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_12e08f07),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_620ff4d8[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_3b19420 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_620ff4d8[0]),
    .e(al_620ff4d8[1]),
    .f(al_620ff4d8[2]),
    .o(al_f4446f72));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_7bda04fa (
    .a(al_f4446f72),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_620ff4d8[3]),
    .f(al_620ff4d8[4]),
    .o(al_65335fa7));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_93eadb35 (
    .a(al_65335fa7),
    .b(al_620ff4d8[5]),
    .c(al_5b144427),
    .d(al_b2febcce[0]),
    .o(al_df8c0cc2));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_124ee5b8 (
    .a(al_df8c0cc2),
    .b(al_620ff4d8[0]),
    .c(al_620ff4d8[1]),
    .o(al_8e20c85e));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_4c26fdb8 (
    .a(al_8e20c85e),
    .b(al_6db5b9d2),
    .c(al_620ff4d8[2]),
    .d(al_620ff4d8[3]),
    .e(al_620ff4d8[4]),
    .o(al_3e72c22b));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_870f5fd6 (
    .a(al_8e20c85e),
    .b(al_6db5b9d2),
    .c(al_620ff4d8[2]),
    .d(al_620ff4d8[3]),
    .o(al_c958e833));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_48074d57 (
    .a(al_df8c0cc2),
    .b(al_6db5b9d2),
    .c(al_620ff4d8[0]),
    .o(al_65670e55));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_1213c38 (
    .a(al_df8c0cc2),
    .b(al_6db5b9d2),
    .c(al_620ff4d8[0]),
    .d(al_620ff4d8[1]),
    .o(al_15ca3484));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_7fe8b7d3 (
    .a(al_8e20c85e),
    .b(al_6db5b9d2),
    .c(al_620ff4d8[2]),
    .o(al_e49c184e));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_918bda78 (
    .a(al_8e20c85e),
    .b(al_6db5b9d2),
    .c(al_620ff4d8[2]),
    .d(al_620ff4d8[3]),
    .e(al_620ff4d8[4]),
    .f(al_620ff4d8[5]),
    .o(al_12e08f07));
  AL_DFF_0 al_b597a472 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_65670e55),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_620ff4d8[0]));
  AL_DFF_0 al_f002d1ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_15ca3484),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_620ff4d8[1]));
  AL_DFF_0 al_aaa68615 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e531b722),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8e42692a[2]));
  AL_DFF_0 al_68b59fe2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e8ea4a8d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8e42692a[3]));
  AL_DFF_0 al_37c2f338 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7d8911c3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8e42692a[4]));
  AL_DFF_0 al_ba8d0064 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4ebe4f9a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d62bafb2[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_a410cdba (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_8e42692a[0]),
    .e(al_8e42692a[1]),
    .f(al_8e42692a[2]),
    .o(al_9c945a81));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_b0f21aab (
    .a(al_9c945a81),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_8e42692a[3]),
    .f(al_8e42692a[4]),
    .o(al_a8eab0c8));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_a28afb01 (
    .a(al_a8eab0c8),
    .b(al_d62bafb2[5]),
    .c(al_42d963e6),
    .d(al_4caca369[0]),
    .o(al_6567b0f6));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_3ddea713 (
    .a(al_6567b0f6),
    .b(al_8e42692a[0]),
    .c(al_8e42692a[1]),
    .d(al_8e42692a[2]),
    .e(al_8e42692a[3]),
    .f(al_8e42692a[4]),
    .o(al_72329cb5));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_66453876 (
    .a(al_6567b0f6),
    .b(al_8e42692a[0]),
    .c(al_8e42692a[1]),
    .d(al_8e42692a[2]),
    .e(al_8e42692a[3]),
    .f(al_8e42692a[4]),
    .o(al_2f10c83f));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_385a70e1 (
    .a(al_2f10c83f),
    .b(al_6db5b9d2),
    .o(al_7d8911c3));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_fdfd5d50 (
    .a(al_6567b0f6),
    .b(al_6db5b9d2),
    .c(al_8e42692a[0]),
    .d(al_8e42692a[1]),
    .e(al_8e42692a[2]),
    .f(al_8e42692a[3]),
    .o(al_e8ea4a8d));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_4fd0c5e5 (
    .a(al_6567b0f6),
    .b(al_6db5b9d2),
    .c(al_8e42692a[0]),
    .o(al_f9924877));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_bf101fc3 (
    .a(al_6567b0f6),
    .b(al_6db5b9d2),
    .c(al_8e42692a[0]),
    .d(al_8e42692a[1]),
    .o(al_26d08bda));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_2b212b64 (
    .a(al_6567b0f6),
    .b(al_6db5b9d2),
    .c(al_8e42692a[0]),
    .d(al_8e42692a[1]),
    .e(al_8e42692a[2]),
    .o(al_e531b722));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_81ed1f67 (
    .a(al_72329cb5),
    .b(al_6db5b9d2),
    .c(al_d62bafb2[5]),
    .o(al_4ebe4f9a));
  AL_DFF_0 al_b948106f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f9924877),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8e42692a[0]));
  AL_DFF_0 al_7f5f5ff7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_26d08bda),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8e42692a[1]));
  AL_DFF_0 al_19577cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_177e297a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5362aaf[2]));
  AL_DFF_0 al_48d33c58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_14d0a20a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5362aaf[3]));
  AL_DFF_0 al_732837aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a855268a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5362aaf[4]));
  AL_DFF_0 al_ee59c07b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4476a641),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5362aaf[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_fd9684b (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_5362aaf[0]),
    .e(al_5362aaf[1]),
    .f(al_5362aaf[2]),
    .o(al_5de748fa));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_6acfccaa (
    .a(al_5de748fa),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_5362aaf[3]),
    .f(al_5362aaf[4]),
    .o(al_d2cdc7c9));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_f18254ac (
    .a(al_d2cdc7c9),
    .b(al_5362aaf[5]),
    .c(al_9a6187ef),
    .d(al_4caca369[0]),
    .o(al_33a1ab04));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_f471a458 (
    .a(al_33a1ab04),
    .b(al_5362aaf[0]),
    .c(al_5362aaf[1]),
    .o(al_ebd8858));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_2e5f775e (
    .a(al_ebd8858),
    .b(al_6db5b9d2),
    .c(al_5362aaf[2]),
    .d(al_5362aaf[3]),
    .e(al_5362aaf[4]),
    .o(al_a855268a));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_74134f8d (
    .a(al_ebd8858),
    .b(al_6db5b9d2),
    .c(al_5362aaf[2]),
    .d(al_5362aaf[3]),
    .o(al_14d0a20a));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_3dd92d3f (
    .a(al_33a1ab04),
    .b(al_6db5b9d2),
    .c(al_5362aaf[0]),
    .o(al_e250e193));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_cdf587b6 (
    .a(al_33a1ab04),
    .b(al_6db5b9d2),
    .c(al_5362aaf[0]),
    .d(al_5362aaf[1]),
    .o(al_c4db602d));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_b7caffba (
    .a(al_ebd8858),
    .b(al_6db5b9d2),
    .c(al_5362aaf[2]),
    .o(al_177e297a));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_6479ce1c (
    .a(al_ebd8858),
    .b(al_6db5b9d2),
    .c(al_5362aaf[2]),
    .d(al_5362aaf[3]),
    .e(al_5362aaf[4]),
    .f(al_5362aaf[5]),
    .o(al_4476a641));
  AL_DFF_0 al_cd0024a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e250e193),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5362aaf[0]));
  AL_DFF_0 al_317931ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c4db602d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5362aaf[1]));
  AL_DFF_0 al_5195a3a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_bb7bf12),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_880139ce[2]));
  AL_DFF_0 al_13d783b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1e407f5a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_880139ce[3]));
  AL_DFF_0 al_286479fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b57079f2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_880139ce[4]));
  AL_DFF_0 al_b4e48a4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b47584c8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d7eff71[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_797cc65e (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_880139ce[0]),
    .e(al_880139ce[1]),
    .f(al_880139ce[2]),
    .o(al_a2eb56c3));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_44f1ba9e (
    .a(al_a2eb56c3),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_880139ce[3]),
    .f(al_880139ce[4]),
    .o(al_c18c53ba));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_c28621e2 (
    .a(al_c18c53ba),
    .b(al_5d7eff71[5]),
    .c(al_f1015bac),
    .d(al_b065182c[0]),
    .o(al_68105619));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_fdaf4d5c (
    .a(al_68105619),
    .b(al_880139ce[0]),
    .c(al_880139ce[1]),
    .o(al_386fccc3));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_62ca269f (
    .a(al_386fccc3),
    .b(al_6db5b9d2),
    .c(al_880139ce[2]),
    .d(al_880139ce[3]),
    .e(al_880139ce[4]),
    .o(al_b57079f2));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_1d535e65 (
    .a(al_386fccc3),
    .b(al_6db5b9d2),
    .c(al_880139ce[2]),
    .d(al_880139ce[3]),
    .o(al_1e407f5a));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_b963d642 (
    .a(al_68105619),
    .b(al_6db5b9d2),
    .c(al_880139ce[0]),
    .o(al_f34da80b));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_3bb26bf2 (
    .a(al_68105619),
    .b(al_6db5b9d2),
    .c(al_880139ce[0]),
    .d(al_880139ce[1]),
    .o(al_df31c3a1));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_d3ba9641 (
    .a(al_386fccc3),
    .b(al_6db5b9d2),
    .c(al_880139ce[2]),
    .o(al_bb7bf12));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_a1dfcd3 (
    .a(al_386fccc3),
    .b(al_6db5b9d2),
    .c(al_880139ce[2]),
    .d(al_880139ce[3]),
    .e(al_880139ce[4]),
    .f(al_5d7eff71[5]),
    .o(al_b47584c8));
  AL_DFF_0 al_3a684178 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f34da80b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_880139ce[0]));
  AL_DFF_0 al_8ca13fdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_df31c3a1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_880139ce[1]));
  AL_DFF_0 al_9051d2a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_53cc0ecc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8119a127[2]));
  AL_DFF_0 al_48354b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2ca2d7bc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8119a127[3]));
  AL_DFF_0 al_42d6fe2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f7fcf2a1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8119a127[4]));
  AL_DFF_0 al_49a7b946 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fdb8587d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd20e4f2[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_34ac5922 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_8119a127[0]),
    .e(al_8119a127[1]),
    .f(al_8119a127[2]),
    .o(al_fb87711d));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_f5eb3239 (
    .a(al_fb87711d),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_8119a127[3]),
    .f(al_8119a127[4]),
    .o(al_38452a92));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_ca853e03 (
    .a(al_38452a92),
    .b(al_dd20e4f2[5]),
    .c(al_8cf002a4),
    .d(al_28515a17[0]),
    .o(al_b0b78459));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_4941b7df (
    .a(al_b0b78459),
    .b(al_8119a127[0]),
    .c(al_8119a127[1]),
    .o(al_6c84cbad));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_11bc6ce1 (
    .a(al_6c84cbad),
    .b(al_6db5b9d2),
    .c(al_8119a127[2]),
    .d(al_8119a127[3]),
    .e(al_8119a127[4]),
    .o(al_f7fcf2a1));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_cf22a4a4 (
    .a(al_6c84cbad),
    .b(al_6db5b9d2),
    .c(al_8119a127[2]),
    .d(al_8119a127[3]),
    .o(al_2ca2d7bc));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_a5f39225 (
    .a(al_b0b78459),
    .b(al_6db5b9d2),
    .c(al_8119a127[0]),
    .o(al_cc8bc87f));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_bc320c07 (
    .a(al_b0b78459),
    .b(al_6db5b9d2),
    .c(al_8119a127[0]),
    .d(al_8119a127[1]),
    .o(al_759d9780));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_91cbade5 (
    .a(al_6c84cbad),
    .b(al_6db5b9d2),
    .c(al_8119a127[2]),
    .o(al_53cc0ecc));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_ac0a8ca0 (
    .a(al_6c84cbad),
    .b(al_6db5b9d2),
    .c(al_8119a127[2]),
    .d(al_8119a127[3]),
    .e(al_8119a127[4]),
    .f(al_dd20e4f2[5]),
    .o(al_fdb8587d));
  AL_DFF_0 al_28bd723a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cc8bc87f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8119a127[0]));
  AL_DFF_0 al_9f2da1ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_759d9780),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8119a127[1]));
  AL_DFF_0 al_b0b70149 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b8a226a2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_17e51133[3]));
  AL_DFF_0 al_54a5d353 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1f6dda96),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_17e51133[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_3f3adf9d (
    .a(al_a7c937ec),
    .b(al_17e51133[0]),
    .c(al_17e51133[1]),
    .o(al_ae23d17f));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_40850758 (
    .a(al_ae23d17f),
    .b(al_6db5b9d2),
    .c(al_17e51133[2]),
    .o(al_41afcc92));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_91eadabd (
    .a(al_a7c937ec),
    .b(al_6db5b9d2),
    .c(al_17e51133[0]),
    .o(al_7fa72a5e));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_228fa9d4 (
    .a(al_a7c937ec),
    .b(al_6db5b9d2),
    .c(al_17e51133[0]),
    .d(al_17e51133[1]),
    .o(al_59879e6b));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_ff905a5 (
    .a(al_ae23d17f),
    .b(al_6db5b9d2),
    .c(al_17e51133[2]),
    .d(al_17e51133[3]),
    .o(al_b8a226a2));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_89b7e973 (
    .a(al_ae23d17f),
    .b(al_6db5b9d2),
    .c(al_17e51133[2]),
    .d(al_17e51133[3]),
    .e(al_17e51133[4]),
    .o(al_1f6dda96));
  AL_DFF_0 al_6f2eeeb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7fa72a5e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_17e51133[0]));
  AL_DFF_0 al_25fa131e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_59879e6b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_17e51133[1]));
  AL_DFF_0 al_d4340834 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_41afcc92),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_17e51133[2]));
  AL_DFF_0 al_2fdef1a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2d126bfd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411ed67e));
  AL_DFF_0 al_6aedee17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2d126bfd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b00f7d00));
  AL_DFF_0 al_d11a11b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2d126bfd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1342f12a));
  AL_DFF_0 al_9ac36373 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c49eb0a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_20e796af));
  AL_DFF_0 al_8baee91c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c49eb0a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f567595c));
  AL_DFF_0 al_105ebdd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c49eb0a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a2b915e0));
  AL_DFF_0 al_24294416 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c49eb0a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d0805f59));
  AL_DFF_0 al_d4f46412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7c49eb0a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_710215be));
  AL_DFF_0 al_27de51a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d6d3de1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5f044880));
  AL_DFF_0 al_ce9d7988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d6d3de1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6e8c75));
  AL_DFF_0 al_c5e692cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d6d3de1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d7411c1e));
  AL_DFF_0 al_93995780 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d6d3de1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dade993));
  AL_DFF_0 al_46f7910b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d6d3de1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ea20fda));
  AL_DFF_0 al_cd50bf0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_151512a8[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9683b2fb));
  AL_DFF_0 al_b830c502 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_151512a8[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e6b3b5a));
  AL_DFF_0 al_49f4e045 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_151512a8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b3b929ae));
  AL_DFF_0 al_f35319f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_151512a8[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb65ad25));
  AL_DFF_0 al_47cfe515 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_151512a8[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_881adcbc));
  AL_DFF_0 al_365b6db5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d23802b0[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_581e4e41[3]));
  AL_DFF_0 al_294e32db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d23802b0[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_581e4e41[4]));
  AL_DFF_0 al_6c697d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d23802b0[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_581e4e41[0]));
  AL_DFF_0 al_57617a77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d23802b0[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_581e4e41[1]));
  AL_DFF_0 al_c1550840 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d23802b0[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_581e4e41[2]));
  AL_DFF_0 al_8b64f6ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_efb91504),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac2df9bf));
  AL_DFF_0 al_97f74bcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_60238e88),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb90ce6));
  AL_DFF_0 al_8c54eae6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_37606c32),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_607ca590));
  AL_DFF_0 al_4b8cb042 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2404250b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33994c72));
  AL_DFF_0 al_f5aaa2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_23e60859),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5082a19[2]));
  AL_DFF_0 al_c7477b91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9cb07372),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5082a19[3]));
  AL_DFF_0 al_6335f74a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cb712978),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5082a19[4]));
  AL_DFF_0 al_8ffea70f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7d870001),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5082a19[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_f81de1fa (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_b5082a19[0]),
    .e(al_b5082a19[1]),
    .f(al_b5082a19[2]),
    .o(al_c254d68a));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_f988cef5 (
    .a(al_c254d68a),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_b5082a19[3]),
    .f(al_b5082a19[4]),
    .o(al_2eb834f5));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_556bd4c6 (
    .a(al_2eb834f5),
    .b(al_b5082a19[5]),
    .c(al_815c8034),
    .d(al_b065182c[0]),
    .o(al_e748e446));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_cd8c4618 (
    .a(al_e748e446),
    .b(al_b5082a19[0]),
    .c(al_b5082a19[1]),
    .o(al_cab235ff));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_ee350b52 (
    .a(al_cab235ff),
    .b(al_6db5b9d2),
    .c(al_b5082a19[2]),
    .d(al_b5082a19[3]),
    .e(al_b5082a19[4]),
    .o(al_cb712978));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_26c6e2fc (
    .a(al_cab235ff),
    .b(al_6db5b9d2),
    .c(al_b5082a19[2]),
    .d(al_b5082a19[3]),
    .o(al_9cb07372));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_ce1daf16 (
    .a(al_e748e446),
    .b(al_6db5b9d2),
    .c(al_b5082a19[0]),
    .o(al_c4e45821));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_3778b44c (
    .a(al_e748e446),
    .b(al_6db5b9d2),
    .c(al_b5082a19[0]),
    .d(al_b5082a19[1]),
    .o(al_aaeb19f7));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_ea7f4d73 (
    .a(al_cab235ff),
    .b(al_6db5b9d2),
    .c(al_b5082a19[2]),
    .o(al_23e60859));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_8e5a3e7b (
    .a(al_cab235ff),
    .b(al_6db5b9d2),
    .c(al_b5082a19[2]),
    .d(al_b5082a19[3]),
    .e(al_b5082a19[4]),
    .f(al_b5082a19[5]),
    .o(al_7d870001));
  AL_DFF_0 al_d2a428eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c4e45821),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5082a19[0]));
  AL_DFF_0 al_dc1cf612 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aaeb19f7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5082a19[1]));
  AL_DFF_0 al_5b423081 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c1ef4c7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a28bab3a));
  AL_DFF_0 al_42dfe7f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_817a8c80),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e0914439));
  AL_DFF_0 al_52c625ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_7e4e201e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_19e026e1[0]));
  AL_DFF_0 al_1f687af0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5b144427),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_19e026e1[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_60edb4ea (
    .a(al_5b144427),
    .b(al_1719553b[0]),
    .o(al_7e4e201e));
  AL_DFF_0 al_80923f5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9681ccaa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48ead91e));
  AL_DFF_0 al_61c400e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1aa44e47[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a390ad74));
  AL_DFF_0 al_3e8b36a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f62892[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c8ccef5));
  AL_DFF_0 al_2f9c1022 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_50ec922d[0]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_41c5883));
  AL_DFF_0 al_3968a6e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_50ec922d[1]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_361b3557));
  AL_DFF_0 al_41f1211e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_50ec922d[2]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_54a8a910));
  AL_DFF_0 al_cb52d75f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_50ec922d[3]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_5f0a94fd));
  AL_DFF_0 al_69ce9b9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_50ec922d[4]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_aa906eb4));
  AL_DFF_0 al_d0f405f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_50ec922d[5]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_20745547));
  AL_DFF_0 al_e6c3d08e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_50ec922d[6]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_8f0f91a1));
  AL_DFF_0 al_c0c33b36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_50ec922d[7]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7d364519));
  AL_DFF_0 al_a3ac80a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d6e96525),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_162fb89b[2]));
  AL_DFF_0 al_1cbbbc6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_224cbb04),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_162fb89b[3]));
  AL_DFF_0 al_ea9ad684 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5c961523),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_162fb89b[4]));
  AL_DFF_0 al_458c1cea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_146bb661),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_162fb89b[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_7fbb2b18 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_162fb89b[0]),
    .e(al_162fb89b[1]),
    .f(al_162fb89b[2]),
    .o(al_ae305841));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_a42a9231 (
    .a(al_ae305841),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_162fb89b[3]),
    .f(al_162fb89b[4]),
    .o(al_a56ffae1));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_b6a9efc8 (
    .a(al_a56ffae1),
    .b(al_162fb89b[5]),
    .c(al_b2febcce[0]),
    .o(al_f5b95ad4));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_ae3d16b3 (
    .a(al_f5b95ad4),
    .b(al_72bfbb1a),
    .o(al_19de37d3));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_ada466f4 (
    .a(al_19de37d3),
    .b(al_162fb89b[0]),
    .c(al_162fb89b[1]),
    .d(al_162fb89b[2]),
    .e(al_162fb89b[3]),
    .f(al_162fb89b[4]),
    .o(al_7b57cbb6));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_8463f8a2 (
    .a(al_19de37d3),
    .b(al_162fb89b[0]),
    .c(al_162fb89b[1]),
    .d(al_162fb89b[2]),
    .e(al_162fb89b[3]),
    .f(al_162fb89b[4]),
    .o(al_b5f76101));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_3e9a528f (
    .a(al_b5f76101),
    .b(al_6db5b9d2),
    .o(al_5c961523));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_f12d7eec (
    .a(al_19de37d3),
    .b(al_6db5b9d2),
    .c(al_162fb89b[0]),
    .d(al_162fb89b[1]),
    .e(al_162fb89b[2]),
    .f(al_162fb89b[3]),
    .o(al_224cbb04));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_2ffb53c2 (
    .a(al_19de37d3),
    .b(al_6db5b9d2),
    .c(al_162fb89b[0]),
    .o(al_a71f7b3c));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_78e1b970 (
    .a(al_19de37d3),
    .b(al_6db5b9d2),
    .c(al_162fb89b[0]),
    .d(al_162fb89b[1]),
    .o(al_6b47e31e));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_d30c588b (
    .a(al_19de37d3),
    .b(al_6db5b9d2),
    .c(al_162fb89b[0]),
    .d(al_162fb89b[1]),
    .e(al_162fb89b[2]),
    .o(al_d6e96525));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_dd72d7ce (
    .a(al_7b57cbb6),
    .b(al_6db5b9d2),
    .c(al_162fb89b[5]),
    .o(al_146bb661));
  AL_DFF_0 al_264d1902 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a71f7b3c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_162fb89b[0]));
  AL_DFF_0 al_69943264 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6b47e31e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_162fb89b[1]));
  AL_DFF_0 al_5085483c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3ca382aa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6b9e41[2]));
  AL_DFF_0 al_99a276a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e5156e61),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6b9e41[3]));
  AL_DFF_0 al_ab2ba56d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_73a263d4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6b9e41[4]));
  AL_DFF_0 al_9bda02de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a502ee6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6b9e41[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_ab935bce (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_d6b9e41[0]),
    .e(al_d6b9e41[1]),
    .f(al_d6b9e41[2]),
    .o(al_73668eea));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_d8e9023e (
    .a(al_73668eea),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_d6b9e41[3]),
    .f(al_d6b9e41[4]),
    .o(al_e3e65c55));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_165cfcf1 (
    .a(al_e3e65c55),
    .b(al_d6b9e41[5]),
    .c(al_87f40037),
    .d(al_28515a17[0]),
    .o(al_6e5fe692));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*~A)"),
    .INIT(64'h4000000000000000))
    al_9a073577 (
    .a(al_6e5fe692),
    .b(al_d6b9e41[0]),
    .c(al_d6b9e41[1]),
    .d(al_d6b9e41[2]),
    .e(al_d6b9e41[3]),
    .f(al_d6b9e41[4]),
    .o(al_9fadbc99));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_e16fff9f (
    .a(al_6e5fe692),
    .b(al_d6b9e41[0]),
    .c(al_d6b9e41[1]),
    .d(al_d6b9e41[2]),
    .e(al_d6b9e41[3]),
    .f(al_d6b9e41[4]),
    .o(al_86543e7b));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_d85aa20f (
    .a(al_86543e7b),
    .b(al_6db5b9d2),
    .o(al_73a263d4));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*~A)))"),
    .INIT(64'h2333333310000000))
    al_eda0e364 (
    .a(al_6e5fe692),
    .b(al_6db5b9d2),
    .c(al_d6b9e41[0]),
    .d(al_d6b9e41[1]),
    .e(al_d6b9e41[2]),
    .f(al_d6b9e41[3]),
    .o(al_e5156e61));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_afd84f77 (
    .a(al_6e5fe692),
    .b(al_6db5b9d2),
    .c(al_d6b9e41[0]),
    .o(al_2c034ec4));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_3a64ef0f (
    .a(al_6e5fe692),
    .b(al_6db5b9d2),
    .c(al_d6b9e41[0]),
    .d(al_d6b9e41[1]),
    .o(al_69054c50));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*~A)))"),
    .INIT(32'h23331000))
    al_58767858 (
    .a(al_6e5fe692),
    .b(al_6db5b9d2),
    .c(al_d6b9e41[0]),
    .d(al_d6b9e41[1]),
    .e(al_d6b9e41[2]),
    .o(al_3ca382aa));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_3aa2dbf4 (
    .a(al_9fadbc99),
    .b(al_6db5b9d2),
    .c(al_d6b9e41[5]),
    .o(al_a502ee6));
  AL_DFF_0 al_668647c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_2c034ec4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6b9e41[0]));
  AL_DFF_0 al_2e6b9de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_69054c50),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6b9e41[1]));
  AL_DFF_0 al_b0a2e05f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_12ccb57b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4206b0c2[2]));
  AL_DFF_0 al_84335f27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4e3c3c1e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4206b0c2[3]));
  AL_DFF_0 al_a62548df (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a68c8fdd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4206b0c2[4]));
  AL_DFF_0 al_639351e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_c6b7617c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4206b0c2[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_3d2149b7 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_4206b0c2[0]),
    .e(al_4206b0c2[1]),
    .f(al_4206b0c2[2]),
    .o(al_ce09b21b));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_4fc0cd10 (
    .a(al_ce09b21b),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_4206b0c2[3]),
    .f(al_4206b0c2[4]),
    .o(al_2c66a236));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_b8ea0db1 (
    .a(al_2c66a236),
    .b(al_4206b0c2[5]),
    .c(al_843f6bac),
    .d(al_4caca369[0]),
    .o(al_7ee2af8f));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_d342e3da (
    .a(al_7ee2af8f),
    .b(al_4206b0c2[0]),
    .c(al_4206b0c2[1]),
    .o(al_10d4c4b6));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_2730f185 (
    .a(al_10d4c4b6),
    .b(al_6db5b9d2),
    .c(al_4206b0c2[2]),
    .d(al_4206b0c2[3]),
    .e(al_4206b0c2[4]),
    .o(al_a68c8fdd));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_8e651026 (
    .a(al_10d4c4b6),
    .b(al_6db5b9d2),
    .c(al_4206b0c2[2]),
    .d(al_4206b0c2[3]),
    .o(al_4e3c3c1e));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_d096ae1f (
    .a(al_7ee2af8f),
    .b(al_6db5b9d2),
    .c(al_4206b0c2[0]),
    .o(al_4d3e12f0));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_26a3d8fd (
    .a(al_7ee2af8f),
    .b(al_6db5b9d2),
    .c(al_4206b0c2[0]),
    .d(al_4206b0c2[1]),
    .o(al_417e5201));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_6d644758 (
    .a(al_10d4c4b6),
    .b(al_6db5b9d2),
    .c(al_4206b0c2[2]),
    .o(al_12ccb57b));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_7bbbbadc (
    .a(al_10d4c4b6),
    .b(al_6db5b9d2),
    .c(al_4206b0c2[2]),
    .d(al_4206b0c2[3]),
    .e(al_4206b0c2[4]),
    .f(al_4206b0c2[5]),
    .o(al_c6b7617c));
  AL_DFF_0 al_6a840016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_4d3e12f0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4206b0c2[0]));
  AL_DFF_0 al_a1da3701 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_417e5201),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4206b0c2[1]));
  AL_DFF_0 al_52e1864a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_94e27914),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44864e28[2]));
  AL_DFF_0 al_2681d730 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8abb9d02),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44864e28[3]));
  AL_DFF_0 al_fbf6ee69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_420e50cb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44864e28[4]));
  AL_DFF_0 al_48bee62b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_42f3bac7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44864e28[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_f050c627 (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_44864e28[0]),
    .e(al_44864e28[1]),
    .f(al_44864e28[2]),
    .o(al_e059f386));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_722f1bdf (
    .a(al_e059f386),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_44864e28[3]),
    .f(al_44864e28[4]),
    .o(al_72450658));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_5d4b7de (
    .a(al_72450658),
    .b(al_44864e28[5]),
    .c(al_535f72cd),
    .d(al_b065182c[0]),
    .o(al_e1983c08));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_54dd5e57 (
    .a(al_e1983c08),
    .b(al_44864e28[0]),
    .c(al_44864e28[1]),
    .o(al_a657a302));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_f185e1dc (
    .a(al_a657a302),
    .b(al_6db5b9d2),
    .c(al_44864e28[2]),
    .d(al_44864e28[3]),
    .e(al_44864e28[4]),
    .o(al_420e50cb));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_5facd206 (
    .a(al_a657a302),
    .b(al_6db5b9d2),
    .c(al_44864e28[2]),
    .d(al_44864e28[3]),
    .o(al_8abb9d02));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_f924930b (
    .a(al_e1983c08),
    .b(al_6db5b9d2),
    .c(al_44864e28[0]),
    .o(al_aefa880a));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_10f2234e (
    .a(al_e1983c08),
    .b(al_6db5b9d2),
    .c(al_44864e28[0]),
    .d(al_44864e28[1]),
    .o(al_dbb207a));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_7d492732 (
    .a(al_a657a302),
    .b(al_6db5b9d2),
    .c(al_44864e28[2]),
    .o(al_94e27914));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_c3cf4d27 (
    .a(al_a657a302),
    .b(al_6db5b9d2),
    .c(al_44864e28[2]),
    .d(al_44864e28[3]),
    .e(al_44864e28[4]),
    .f(al_44864e28[5]),
    .o(al_42f3bac7));
  AL_DFF_0 al_acdbe3fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aefa880a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44864e28[0]));
  AL_DFF_0 al_44a40bc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_dbb207a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44864e28[1]));
  AL_DFF_0 al_1c73acb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9aed2757),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71242bdd[2]));
  AL_DFF_0 al_cd5791ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_ed505fc9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71242bdd[3]));
  AL_DFF_0 al_68acce42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d3c1dd73),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71242bdd[4]));
  AL_DFF_0 al_e6617d8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b76e4bca),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71242bdd[5]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_148352ce (
    .a(al_9841dcd3),
    .b(al_7a04bdba),
    .o(al_99c75e01));
  AL_MAP_LUT6 #(
    .EQN("~(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h7fbfdfeff7fbfdfe))
    al_e0c2a0ec (
    .a(al_511af127[0]),
    .b(al_511af127[1]),
    .c(al_511af127[2]),
    .d(al_71242bdd[0]),
    .e(al_71242bdd[1]),
    .f(al_71242bdd[2]),
    .o(al_31a7d949));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_9b0f36d2 (
    .a(al_31a7d949),
    .b(al_99c75e01),
    .c(al_511af127[3]),
    .d(al_511af127[4]),
    .e(al_71242bdd[3]),
    .f(al_71242bdd[4]),
    .o(al_fd1400b6));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*(D@B))"),
    .INIT(16'h1040))
    al_bc3eff76 (
    .a(al_fd1400b6),
    .b(al_71242bdd[5]),
    .c(al_17b42586),
    .d(al_28515a17[0]),
    .o(al_38d9fe9));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_96516a41 (
    .a(al_38d9fe9),
    .b(al_71242bdd[0]),
    .c(al_71242bdd[1]),
    .o(al_bd9a895c));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_fcf97ab (
    .a(al_bd9a895c),
    .b(al_6db5b9d2),
    .c(al_71242bdd[2]),
    .d(al_71242bdd[3]),
    .e(al_71242bdd[4]),
    .o(al_d3c1dd73));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_1b114695 (
    .a(al_bd9a895c),
    .b(al_6db5b9d2),
    .c(al_71242bdd[2]),
    .d(al_71242bdd[3]),
    .o(al_ed505fc9));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_1db1edf7 (
    .a(al_38d9fe9),
    .b(al_6db5b9d2),
    .c(al_71242bdd[0]),
    .o(al_46228dd4));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_eda22860 (
    .a(al_38d9fe9),
    .b(al_6db5b9d2),
    .c(al_71242bdd[0]),
    .d(al_71242bdd[1]),
    .o(al_d9253b60));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_633749bc (
    .a(al_bd9a895c),
    .b(al_6db5b9d2),
    .c(al_71242bdd[2]),
    .o(al_9aed2757));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_bb9052be (
    .a(al_bd9a895c),
    .b(al_6db5b9d2),
    .c(al_71242bdd[2]),
    .d(al_71242bdd[3]),
    .e(al_71242bdd[4]),
    .f(al_71242bdd[5]),
    .o(al_b76e4bca));
  AL_DFF_0 al_6350af41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_46228dd4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71242bdd[0]));
  AL_DFF_0 al_954fb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d9253b60),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71242bdd[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7af17a28 (
    .a(ddr_app_wdf_data[0]),
    .b(al_8235546f[0]),
    .c(al_e6043332),
    .o(al_c665bb87[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e762dddf (
    .a(ddr_app_wdf_data[100]),
    .b(al_8235546f[100]),
    .c(al_e6043332),
    .o(al_c665bb87[100]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c5ef5592 (
    .a(ddr_app_wdf_data[101]),
    .b(al_8235546f[101]),
    .c(al_e6043332),
    .o(al_c665bb87[101]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e01d6c45 (
    .a(ddr_app_wdf_data[102]),
    .b(al_8235546f[102]),
    .c(al_e6043332),
    .o(al_c665bb87[102]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_75510dbd (
    .a(ddr_app_wdf_data[103]),
    .b(al_8235546f[103]),
    .c(al_e6043332),
    .o(al_c665bb87[103]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e1c61ba8 (
    .a(ddr_app_wdf_data[104]),
    .b(al_8235546f[104]),
    .c(al_e6043332),
    .o(al_c665bb87[104]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8ce5dd15 (
    .a(ddr_app_wdf_data[105]),
    .b(al_8235546f[105]),
    .c(al_e6043332),
    .o(al_c665bb87[105]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_56f14437 (
    .a(ddr_app_wdf_data[106]),
    .b(al_8235546f[106]),
    .c(al_e6043332),
    .o(al_c665bb87[106]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_71812e66 (
    .a(ddr_app_wdf_data[107]),
    .b(al_8235546f[107]),
    .c(al_e6043332),
    .o(al_c665bb87[107]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_beca01b7 (
    .a(ddr_app_wdf_data[108]),
    .b(al_8235546f[108]),
    .c(al_e6043332),
    .o(al_c665bb87[108]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_eb706717 (
    .a(ddr_app_wdf_data[109]),
    .b(al_8235546f[109]),
    .c(al_e6043332),
    .o(al_c665bb87[109]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8786256c (
    .a(ddr_app_wdf_data[10]),
    .b(al_8235546f[10]),
    .c(al_e6043332),
    .o(al_c665bb87[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_266a0d7f (
    .a(ddr_app_wdf_data[110]),
    .b(al_8235546f[110]),
    .c(al_e6043332),
    .o(al_c665bb87[110]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ea6326f4 (
    .a(ddr_app_wdf_data[111]),
    .b(al_8235546f[111]),
    .c(al_e6043332),
    .o(al_c665bb87[111]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3b6c6420 (
    .a(ddr_app_wdf_data[112]),
    .b(al_8235546f[112]),
    .c(al_e6043332),
    .o(al_c665bb87[112]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d8548da7 (
    .a(ddr_app_wdf_data[113]),
    .b(al_8235546f[113]),
    .c(al_e6043332),
    .o(al_c665bb87[113]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_dbc742c1 (
    .a(ddr_app_wdf_data[114]),
    .b(al_8235546f[114]),
    .c(al_e6043332),
    .o(al_c665bb87[114]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_87cc4e90 (
    .a(ddr_app_wdf_data[115]),
    .b(al_8235546f[115]),
    .c(al_e6043332),
    .o(al_c665bb87[115]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8254019 (
    .a(ddr_app_wdf_data[116]),
    .b(al_8235546f[116]),
    .c(al_e6043332),
    .o(al_c665bb87[116]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a0d2a134 (
    .a(ddr_app_wdf_data[117]),
    .b(al_8235546f[117]),
    .c(al_e6043332),
    .o(al_c665bb87[117]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e5852b71 (
    .a(ddr_app_wdf_data[118]),
    .b(al_8235546f[118]),
    .c(al_e6043332),
    .o(al_c665bb87[118]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c9ff313 (
    .a(ddr_app_wdf_data[119]),
    .b(al_8235546f[119]),
    .c(al_e6043332),
    .o(al_c665bb87[119]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ffcb179b (
    .a(ddr_app_wdf_data[11]),
    .b(al_8235546f[11]),
    .c(al_e6043332),
    .o(al_c665bb87[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_47283fa3 (
    .a(ddr_app_wdf_data[120]),
    .b(al_8235546f[120]),
    .c(al_e6043332),
    .o(al_c665bb87[120]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_331900c8 (
    .a(ddr_app_wdf_data[121]),
    .b(al_8235546f[121]),
    .c(al_e6043332),
    .o(al_c665bb87[121]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d0e03d4 (
    .a(ddr_app_wdf_data[122]),
    .b(al_8235546f[122]),
    .c(al_e6043332),
    .o(al_c665bb87[122]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e088cff8 (
    .a(ddr_app_wdf_data[123]),
    .b(al_8235546f[123]),
    .c(al_e6043332),
    .o(al_c665bb87[123]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_bb7605fb (
    .a(ddr_app_wdf_data[124]),
    .b(al_8235546f[124]),
    .c(al_e6043332),
    .o(al_c665bb87[124]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a875d7fa (
    .a(ddr_app_wdf_data[125]),
    .b(al_8235546f[125]),
    .c(al_e6043332),
    .o(al_c665bb87[125]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e789059e (
    .a(ddr_app_wdf_data[126]),
    .b(al_8235546f[126]),
    .c(al_e6043332),
    .o(al_c665bb87[126]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f3814de7 (
    .a(ddr_app_wdf_data[127]),
    .b(al_8235546f[127]),
    .c(al_e6043332),
    .o(al_c665bb87[127]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fc4e3361 (
    .a(ddr_app_wdf_data[128]),
    .b(al_8235546f[128]),
    .c(al_e6043332),
    .o(al_c665bb87[128]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3f50d39f (
    .a(ddr_app_wdf_data[129]),
    .b(al_8235546f[129]),
    .c(al_e6043332),
    .o(al_c665bb87[129]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3c2d30e6 (
    .a(ddr_app_wdf_data[12]),
    .b(al_8235546f[12]),
    .c(al_e6043332),
    .o(al_c665bb87[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b5c1bd6a (
    .a(ddr_app_wdf_data[130]),
    .b(al_8235546f[130]),
    .c(al_e6043332),
    .o(al_c665bb87[130]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e40c34e6 (
    .a(ddr_app_wdf_data[131]),
    .b(al_8235546f[131]),
    .c(al_e6043332),
    .o(al_c665bb87[131]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7bcc52e7 (
    .a(ddr_app_wdf_data[132]),
    .b(al_8235546f[132]),
    .c(al_e6043332),
    .o(al_c665bb87[132]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e0e4e057 (
    .a(ddr_app_wdf_data[133]),
    .b(al_8235546f[133]),
    .c(al_e6043332),
    .o(al_c665bb87[133]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2a4ee126 (
    .a(ddr_app_wdf_data[134]),
    .b(al_8235546f[134]),
    .c(al_e6043332),
    .o(al_c665bb87[134]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4d98a7ff (
    .a(ddr_app_wdf_data[135]),
    .b(al_8235546f[135]),
    .c(al_e6043332),
    .o(al_c665bb87[135]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1c6d20f0 (
    .a(ddr_app_wdf_data[136]),
    .b(al_8235546f[136]),
    .c(al_e6043332),
    .o(al_c665bb87[136]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_17981b67 (
    .a(ddr_app_wdf_data[137]),
    .b(al_8235546f[137]),
    .c(al_e6043332),
    .o(al_c665bb87[137]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_944d0716 (
    .a(ddr_app_wdf_data[138]),
    .b(al_8235546f[138]),
    .c(al_e6043332),
    .o(al_c665bb87[138]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1c45fdad (
    .a(ddr_app_wdf_data[139]),
    .b(al_8235546f[139]),
    .c(al_e6043332),
    .o(al_c665bb87[139]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b54153ec (
    .a(ddr_app_wdf_data[13]),
    .b(al_8235546f[13]),
    .c(al_e6043332),
    .o(al_c665bb87[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f8623cfe (
    .a(ddr_app_wdf_data[140]),
    .b(al_8235546f[140]),
    .c(al_e6043332),
    .o(al_c665bb87[140]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_81424f5a (
    .a(ddr_app_wdf_data[141]),
    .b(al_8235546f[141]),
    .c(al_e6043332),
    .o(al_c665bb87[141]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_93b13cd7 (
    .a(ddr_app_wdf_data[142]),
    .b(al_8235546f[142]),
    .c(al_e6043332),
    .o(al_c665bb87[142]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f36d53e2 (
    .a(ddr_app_wdf_data[143]),
    .b(al_8235546f[143]),
    .c(al_e6043332),
    .o(al_c665bb87[143]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d8b38fc (
    .a(ddr_app_wdf_data[144]),
    .b(al_8235546f[144]),
    .c(al_e6043332),
    .o(al_c665bb87[144]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e051171c (
    .a(ddr_app_wdf_data[145]),
    .b(al_8235546f[145]),
    .c(al_e6043332),
    .o(al_c665bb87[145]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f6499203 (
    .a(ddr_app_wdf_data[146]),
    .b(al_8235546f[146]),
    .c(al_e6043332),
    .o(al_c665bb87[146]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_752df8ed (
    .a(ddr_app_wdf_data[147]),
    .b(al_8235546f[147]),
    .c(al_e6043332),
    .o(al_c665bb87[147]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5013a9d6 (
    .a(ddr_app_wdf_data[148]),
    .b(al_8235546f[148]),
    .c(al_e6043332),
    .o(al_c665bb87[148]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c19d8871 (
    .a(ddr_app_wdf_data[149]),
    .b(al_8235546f[149]),
    .c(al_e6043332),
    .o(al_c665bb87[149]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fbf9f1b9 (
    .a(ddr_app_wdf_data[14]),
    .b(al_8235546f[14]),
    .c(al_e6043332),
    .o(al_c665bb87[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7396a443 (
    .a(ddr_app_wdf_data[150]),
    .b(al_8235546f[150]),
    .c(al_e6043332),
    .o(al_c665bb87[150]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ab35b056 (
    .a(ddr_app_wdf_data[151]),
    .b(al_8235546f[151]),
    .c(al_e6043332),
    .o(al_c665bb87[151]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4287c41e (
    .a(ddr_app_wdf_data[152]),
    .b(al_8235546f[152]),
    .c(al_e6043332),
    .o(al_c665bb87[152]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c92976a6 (
    .a(ddr_app_wdf_data[153]),
    .b(al_8235546f[153]),
    .c(al_e6043332),
    .o(al_c665bb87[153]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_93e5b6dc (
    .a(ddr_app_wdf_data[154]),
    .b(al_8235546f[154]),
    .c(al_e6043332),
    .o(al_c665bb87[154]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d5d02ed (
    .a(ddr_app_wdf_data[155]),
    .b(al_8235546f[155]),
    .c(al_e6043332),
    .o(al_c665bb87[155]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_10a251b6 (
    .a(ddr_app_wdf_data[156]),
    .b(al_8235546f[156]),
    .c(al_e6043332),
    .o(al_c665bb87[156]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3789f81d (
    .a(ddr_app_wdf_data[157]),
    .b(al_8235546f[157]),
    .c(al_e6043332),
    .o(al_c665bb87[157]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_19f5f1a4 (
    .a(ddr_app_wdf_data[158]),
    .b(al_8235546f[158]),
    .c(al_e6043332),
    .o(al_c665bb87[158]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c5940895 (
    .a(ddr_app_wdf_data[159]),
    .b(al_8235546f[159]),
    .c(al_e6043332),
    .o(al_c665bb87[159]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a071ba09 (
    .a(ddr_app_wdf_data[15]),
    .b(al_8235546f[15]),
    .c(al_e6043332),
    .o(al_c665bb87[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c61a857b (
    .a(ddr_app_wdf_data[160]),
    .b(al_8235546f[160]),
    .c(al_e6043332),
    .o(al_c665bb87[160]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7b3e07f (
    .a(ddr_app_wdf_data[161]),
    .b(al_8235546f[161]),
    .c(al_e6043332),
    .o(al_c665bb87[161]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c137d095 (
    .a(ddr_app_wdf_data[162]),
    .b(al_8235546f[162]),
    .c(al_e6043332),
    .o(al_c665bb87[162]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_db7def48 (
    .a(ddr_app_wdf_data[163]),
    .b(al_8235546f[163]),
    .c(al_e6043332),
    .o(al_c665bb87[163]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a9527997 (
    .a(ddr_app_wdf_data[164]),
    .b(al_8235546f[164]),
    .c(al_e6043332),
    .o(al_c665bb87[164]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_16e6693c (
    .a(ddr_app_wdf_data[165]),
    .b(al_8235546f[165]),
    .c(al_e6043332),
    .o(al_c665bb87[165]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3e4e35e0 (
    .a(ddr_app_wdf_data[166]),
    .b(al_8235546f[166]),
    .c(al_e6043332),
    .o(al_c665bb87[166]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_cf5e68b9 (
    .a(ddr_app_wdf_data[167]),
    .b(al_8235546f[167]),
    .c(al_e6043332),
    .o(al_c665bb87[167]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3584d427 (
    .a(ddr_app_wdf_data[168]),
    .b(al_8235546f[168]),
    .c(al_e6043332),
    .o(al_c665bb87[168]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_177a8bf5 (
    .a(ddr_app_wdf_data[169]),
    .b(al_8235546f[169]),
    .c(al_e6043332),
    .o(al_c665bb87[169]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9caf839b (
    .a(ddr_app_wdf_data[16]),
    .b(al_8235546f[16]),
    .c(al_e6043332),
    .o(al_c665bb87[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f8a68da9 (
    .a(ddr_app_wdf_data[170]),
    .b(al_8235546f[170]),
    .c(al_e6043332),
    .o(al_c665bb87[170]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_88b2d57e (
    .a(ddr_app_wdf_data[171]),
    .b(al_8235546f[171]),
    .c(al_e6043332),
    .o(al_c665bb87[171]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4e196f69 (
    .a(ddr_app_wdf_data[172]),
    .b(al_8235546f[172]),
    .c(al_e6043332),
    .o(al_c665bb87[172]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fb50a8e7 (
    .a(ddr_app_wdf_data[173]),
    .b(al_8235546f[173]),
    .c(al_e6043332),
    .o(al_c665bb87[173]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_21a00a9b (
    .a(ddr_app_wdf_data[174]),
    .b(al_8235546f[174]),
    .c(al_e6043332),
    .o(al_c665bb87[174]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7a3cb54e (
    .a(ddr_app_wdf_data[175]),
    .b(al_8235546f[175]),
    .c(al_e6043332),
    .o(al_c665bb87[175]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_79be7e02 (
    .a(ddr_app_wdf_data[176]),
    .b(al_8235546f[176]),
    .c(al_e6043332),
    .o(al_c665bb87[176]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f1778e63 (
    .a(ddr_app_wdf_data[177]),
    .b(al_8235546f[177]),
    .c(al_e6043332),
    .o(al_c665bb87[177]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_6a58b456 (
    .a(ddr_app_wdf_data[178]),
    .b(al_8235546f[178]),
    .c(al_e6043332),
    .o(al_c665bb87[178]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c7ee6a1d (
    .a(ddr_app_wdf_data[179]),
    .b(al_8235546f[179]),
    .c(al_e6043332),
    .o(al_c665bb87[179]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7d4a63aa (
    .a(ddr_app_wdf_data[17]),
    .b(al_8235546f[17]),
    .c(al_e6043332),
    .o(al_c665bb87[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ef8f30d (
    .a(ddr_app_wdf_data[180]),
    .b(al_8235546f[180]),
    .c(al_e6043332),
    .o(al_c665bb87[180]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_dbb8b24c (
    .a(ddr_app_wdf_data[181]),
    .b(al_8235546f[181]),
    .c(al_e6043332),
    .o(al_c665bb87[181]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8a583b83 (
    .a(ddr_app_wdf_data[182]),
    .b(al_8235546f[182]),
    .c(al_e6043332),
    .o(al_c665bb87[182]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b562c8d4 (
    .a(ddr_app_wdf_data[183]),
    .b(al_8235546f[183]),
    .c(al_e6043332),
    .o(al_c665bb87[183]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a000615b (
    .a(ddr_app_wdf_data[184]),
    .b(al_8235546f[184]),
    .c(al_e6043332),
    .o(al_c665bb87[184]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f15415d1 (
    .a(ddr_app_wdf_data[185]),
    .b(al_8235546f[185]),
    .c(al_e6043332),
    .o(al_c665bb87[185]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_dd244cc4 (
    .a(ddr_app_wdf_data[186]),
    .b(al_8235546f[186]),
    .c(al_e6043332),
    .o(al_c665bb87[186]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9461e12f (
    .a(ddr_app_wdf_data[187]),
    .b(al_8235546f[187]),
    .c(al_e6043332),
    .o(al_c665bb87[187]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3f10e205 (
    .a(ddr_app_wdf_data[188]),
    .b(al_8235546f[188]),
    .c(al_e6043332),
    .o(al_c665bb87[188]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_57d73208 (
    .a(ddr_app_wdf_data[189]),
    .b(al_8235546f[189]),
    .c(al_e6043332),
    .o(al_c665bb87[189]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_affa2cba (
    .a(ddr_app_wdf_data[18]),
    .b(al_8235546f[18]),
    .c(al_e6043332),
    .o(al_c665bb87[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_904263dd (
    .a(ddr_app_wdf_data[190]),
    .b(al_8235546f[190]),
    .c(al_e6043332),
    .o(al_c665bb87[190]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fc88b16d (
    .a(ddr_app_wdf_data[191]),
    .b(al_8235546f[191]),
    .c(al_e6043332),
    .o(al_c665bb87[191]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3dd88a37 (
    .a(ddr_app_wdf_data[192]),
    .b(al_8235546f[192]),
    .c(al_e6043332),
    .o(al_c665bb87[192]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c014173c (
    .a(ddr_app_wdf_data[193]),
    .b(al_8235546f[193]),
    .c(al_e6043332),
    .o(al_c665bb87[193]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ceea72f5 (
    .a(ddr_app_wdf_data[194]),
    .b(al_8235546f[194]),
    .c(al_e6043332),
    .o(al_c665bb87[194]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_728d5c2b (
    .a(ddr_app_wdf_data[195]),
    .b(al_8235546f[195]),
    .c(al_e6043332),
    .o(al_c665bb87[195]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_20dfc2c1 (
    .a(ddr_app_wdf_data[196]),
    .b(al_8235546f[196]),
    .c(al_e6043332),
    .o(al_c665bb87[196]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_10d14b0a (
    .a(ddr_app_wdf_data[197]),
    .b(al_8235546f[197]),
    .c(al_e6043332),
    .o(al_c665bb87[197]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_dfa04ed6 (
    .a(ddr_app_wdf_data[198]),
    .b(al_8235546f[198]),
    .c(al_e6043332),
    .o(al_c665bb87[198]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_78a0814b (
    .a(ddr_app_wdf_data[199]),
    .b(al_8235546f[199]),
    .c(al_e6043332),
    .o(al_c665bb87[199]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b62551d6 (
    .a(ddr_app_wdf_data[19]),
    .b(al_8235546f[19]),
    .c(al_e6043332),
    .o(al_c665bb87[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c145f1d4 (
    .a(ddr_app_wdf_data[1]),
    .b(al_8235546f[1]),
    .c(al_e6043332),
    .o(al_c665bb87[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d1bd2b98 (
    .a(ddr_app_wdf_data[200]),
    .b(al_8235546f[200]),
    .c(al_e6043332),
    .o(al_c665bb87[200]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_20d5b617 (
    .a(ddr_app_wdf_data[201]),
    .b(al_8235546f[201]),
    .c(al_e6043332),
    .o(al_c665bb87[201]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1f541858 (
    .a(ddr_app_wdf_data[202]),
    .b(al_8235546f[202]),
    .c(al_e6043332),
    .o(al_c665bb87[202]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_69a31ea1 (
    .a(ddr_app_wdf_data[203]),
    .b(al_8235546f[203]),
    .c(al_e6043332),
    .o(al_c665bb87[203]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a86a6945 (
    .a(ddr_app_wdf_data[204]),
    .b(al_8235546f[204]),
    .c(al_e6043332),
    .o(al_c665bb87[204]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7db53540 (
    .a(ddr_app_wdf_data[205]),
    .b(al_8235546f[205]),
    .c(al_e6043332),
    .o(al_c665bb87[205]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d5e2deb3 (
    .a(ddr_app_wdf_data[206]),
    .b(al_8235546f[206]),
    .c(al_e6043332),
    .o(al_c665bb87[206]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4206cee4 (
    .a(ddr_app_wdf_data[207]),
    .b(al_8235546f[207]),
    .c(al_e6043332),
    .o(al_c665bb87[207]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e55bc42c (
    .a(ddr_app_wdf_data[208]),
    .b(al_8235546f[208]),
    .c(al_e6043332),
    .o(al_c665bb87[208]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e140f16d (
    .a(ddr_app_wdf_data[209]),
    .b(al_8235546f[209]),
    .c(al_e6043332),
    .o(al_c665bb87[209]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2d42e200 (
    .a(ddr_app_wdf_data[20]),
    .b(al_8235546f[20]),
    .c(al_e6043332),
    .o(al_c665bb87[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ab1449c9 (
    .a(ddr_app_wdf_data[210]),
    .b(al_8235546f[210]),
    .c(al_e6043332),
    .o(al_c665bb87[210]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1880f18d (
    .a(ddr_app_wdf_data[211]),
    .b(al_8235546f[211]),
    .c(al_e6043332),
    .o(al_c665bb87[211]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_96a462ea (
    .a(ddr_app_wdf_data[212]),
    .b(al_8235546f[212]),
    .c(al_e6043332),
    .o(al_c665bb87[212]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_66005cde (
    .a(ddr_app_wdf_data[213]),
    .b(al_8235546f[213]),
    .c(al_e6043332),
    .o(al_c665bb87[213]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_54cbbd7c (
    .a(ddr_app_wdf_data[214]),
    .b(al_8235546f[214]),
    .c(al_e6043332),
    .o(al_c665bb87[214]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a7995f0f (
    .a(ddr_app_wdf_data[215]),
    .b(al_8235546f[215]),
    .c(al_e6043332),
    .o(al_c665bb87[215]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3f80fa81 (
    .a(ddr_app_wdf_data[216]),
    .b(al_8235546f[216]),
    .c(al_e6043332),
    .o(al_c665bb87[216]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fe94a24b (
    .a(ddr_app_wdf_data[217]),
    .b(al_8235546f[217]),
    .c(al_e6043332),
    .o(al_c665bb87[217]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_88f2f5c0 (
    .a(ddr_app_wdf_data[218]),
    .b(al_8235546f[218]),
    .c(al_e6043332),
    .o(al_c665bb87[218]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7d5f272 (
    .a(ddr_app_wdf_data[219]),
    .b(al_8235546f[219]),
    .c(al_e6043332),
    .o(al_c665bb87[219]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8df06148 (
    .a(ddr_app_wdf_data[21]),
    .b(al_8235546f[21]),
    .c(al_e6043332),
    .o(al_c665bb87[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8533d07d (
    .a(ddr_app_wdf_data[220]),
    .b(al_8235546f[220]),
    .c(al_e6043332),
    .o(al_c665bb87[220]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3892b6b1 (
    .a(ddr_app_wdf_data[221]),
    .b(al_8235546f[221]),
    .c(al_e6043332),
    .o(al_c665bb87[221]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_21131752 (
    .a(ddr_app_wdf_data[222]),
    .b(al_8235546f[222]),
    .c(al_e6043332),
    .o(al_c665bb87[222]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ba557a2d (
    .a(ddr_app_wdf_data[223]),
    .b(al_8235546f[223]),
    .c(al_e6043332),
    .o(al_c665bb87[223]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_eb52dc47 (
    .a(ddr_app_wdf_data[224]),
    .b(al_8235546f[224]),
    .c(al_e6043332),
    .o(al_c665bb87[224]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_40b45e5e (
    .a(ddr_app_wdf_data[225]),
    .b(al_8235546f[225]),
    .c(al_e6043332),
    .o(al_c665bb87[225]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a3f46cc5 (
    .a(ddr_app_wdf_data[226]),
    .b(al_8235546f[226]),
    .c(al_e6043332),
    .o(al_c665bb87[226]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_dcafe3e6 (
    .a(ddr_app_wdf_data[227]),
    .b(al_8235546f[227]),
    .c(al_e6043332),
    .o(al_c665bb87[227]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3b60263e (
    .a(ddr_app_wdf_data[228]),
    .b(al_8235546f[228]),
    .c(al_e6043332),
    .o(al_c665bb87[228]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d4184f07 (
    .a(ddr_app_wdf_data[229]),
    .b(al_8235546f[229]),
    .c(al_e6043332),
    .o(al_c665bb87[229]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2bbdfedc (
    .a(ddr_app_wdf_data[22]),
    .b(al_8235546f[22]),
    .c(al_e6043332),
    .o(al_c665bb87[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9aea894b (
    .a(ddr_app_wdf_data[230]),
    .b(al_8235546f[230]),
    .c(al_e6043332),
    .o(al_c665bb87[230]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a829e383 (
    .a(ddr_app_wdf_data[231]),
    .b(al_8235546f[231]),
    .c(al_e6043332),
    .o(al_c665bb87[231]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8ba4e30a (
    .a(ddr_app_wdf_data[232]),
    .b(al_8235546f[232]),
    .c(al_e6043332),
    .o(al_c665bb87[232]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3261213 (
    .a(ddr_app_wdf_data[233]),
    .b(al_8235546f[233]),
    .c(al_e6043332),
    .o(al_c665bb87[233]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_99d92deb (
    .a(ddr_app_wdf_data[234]),
    .b(al_8235546f[234]),
    .c(al_e6043332),
    .o(al_c665bb87[234]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1674b46e (
    .a(ddr_app_wdf_data[235]),
    .b(al_8235546f[235]),
    .c(al_e6043332),
    .o(al_c665bb87[235]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8ce7f837 (
    .a(ddr_app_wdf_data[236]),
    .b(al_8235546f[236]),
    .c(al_e6043332),
    .o(al_c665bb87[236]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b35d89bf (
    .a(ddr_app_wdf_data[237]),
    .b(al_8235546f[237]),
    .c(al_e6043332),
    .o(al_c665bb87[237]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b74e8075 (
    .a(ddr_app_wdf_data[238]),
    .b(al_8235546f[238]),
    .c(al_e6043332),
    .o(al_c665bb87[238]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f24eec07 (
    .a(ddr_app_wdf_data[239]),
    .b(al_8235546f[239]),
    .c(al_e6043332),
    .o(al_c665bb87[239]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c99b08f6 (
    .a(ddr_app_wdf_data[23]),
    .b(al_8235546f[23]),
    .c(al_e6043332),
    .o(al_c665bb87[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c1f80d56 (
    .a(ddr_app_wdf_data[240]),
    .b(al_8235546f[240]),
    .c(al_e6043332),
    .o(al_c665bb87[240]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_534b56d3 (
    .a(ddr_app_wdf_data[241]),
    .b(al_8235546f[241]),
    .c(al_e6043332),
    .o(al_c665bb87[241]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fea0ba74 (
    .a(ddr_app_wdf_data[242]),
    .b(al_8235546f[242]),
    .c(al_e6043332),
    .o(al_c665bb87[242]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f00fe76 (
    .a(ddr_app_wdf_data[243]),
    .b(al_8235546f[243]),
    .c(al_e6043332),
    .o(al_c665bb87[243]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_6fc5474b (
    .a(ddr_app_wdf_data[244]),
    .b(al_8235546f[244]),
    .c(al_e6043332),
    .o(al_c665bb87[244]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2b70e4fe (
    .a(ddr_app_wdf_data[245]),
    .b(al_8235546f[245]),
    .c(al_e6043332),
    .o(al_c665bb87[245]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7fe0939c (
    .a(ddr_app_wdf_data[246]),
    .b(al_8235546f[246]),
    .c(al_e6043332),
    .o(al_c665bb87[246]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ce7c90f3 (
    .a(ddr_app_wdf_data[247]),
    .b(al_8235546f[247]),
    .c(al_e6043332),
    .o(al_c665bb87[247]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5e5844b7 (
    .a(ddr_app_wdf_data[248]),
    .b(al_8235546f[248]),
    .c(al_e6043332),
    .o(al_c665bb87[248]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_24d180e7 (
    .a(ddr_app_wdf_data[249]),
    .b(al_8235546f[249]),
    .c(al_e6043332),
    .o(al_c665bb87[249]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_caf4a565 (
    .a(ddr_app_wdf_data[24]),
    .b(al_8235546f[24]),
    .c(al_e6043332),
    .o(al_c665bb87[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_818affdc (
    .a(ddr_app_wdf_data[250]),
    .b(al_8235546f[250]),
    .c(al_e6043332),
    .o(al_c665bb87[250]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8cac323d (
    .a(ddr_app_wdf_data[251]),
    .b(al_8235546f[251]),
    .c(al_e6043332),
    .o(al_c665bb87[251]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b62b8749 (
    .a(ddr_app_wdf_data[252]),
    .b(al_8235546f[252]),
    .c(al_e6043332),
    .o(al_c665bb87[252]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_40515e93 (
    .a(ddr_app_wdf_data[253]),
    .b(al_8235546f[253]),
    .c(al_e6043332),
    .o(al_c665bb87[253]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_af496c7d (
    .a(ddr_app_wdf_data[254]),
    .b(al_8235546f[254]),
    .c(al_e6043332),
    .o(al_c665bb87[254]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_99f3065f (
    .a(ddr_app_wdf_data[255]),
    .b(al_8235546f[255]),
    .c(al_e6043332),
    .o(al_c665bb87[255]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_db03d42c (
    .a(ddr_app_wdf_data[25]),
    .b(al_8235546f[25]),
    .c(al_e6043332),
    .o(al_c665bb87[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_230d03e0 (
    .a(ddr_app_wdf_data[26]),
    .b(al_8235546f[26]),
    .c(al_e6043332),
    .o(al_c665bb87[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d6893e2c (
    .a(ddr_app_wdf_data[27]),
    .b(al_8235546f[27]),
    .c(al_e6043332),
    .o(al_c665bb87[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2edd33bf (
    .a(ddr_app_wdf_data[28]),
    .b(al_8235546f[28]),
    .c(al_e6043332),
    .o(al_c665bb87[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_eb7d7d29 (
    .a(ddr_app_wdf_data[29]),
    .b(al_8235546f[29]),
    .c(al_e6043332),
    .o(al_c665bb87[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_73c3124e (
    .a(ddr_app_wdf_data[2]),
    .b(al_8235546f[2]),
    .c(al_e6043332),
    .o(al_c665bb87[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a8e0f793 (
    .a(ddr_app_wdf_data[30]),
    .b(al_8235546f[30]),
    .c(al_e6043332),
    .o(al_c665bb87[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_41cf588d (
    .a(ddr_app_wdf_data[31]),
    .b(al_8235546f[31]),
    .c(al_e6043332),
    .o(al_c665bb87[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1364098d (
    .a(ddr_app_wdf_data[32]),
    .b(al_8235546f[32]),
    .c(al_e6043332),
    .o(al_c665bb87[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_96189a6e (
    .a(ddr_app_wdf_data[33]),
    .b(al_8235546f[33]),
    .c(al_e6043332),
    .o(al_c665bb87[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d37d1181 (
    .a(ddr_app_wdf_data[34]),
    .b(al_8235546f[34]),
    .c(al_e6043332),
    .o(al_c665bb87[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c6ce26aa (
    .a(ddr_app_wdf_data[35]),
    .b(al_8235546f[35]),
    .c(al_e6043332),
    .o(al_c665bb87[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_468fb5f8 (
    .a(ddr_app_wdf_data[36]),
    .b(al_8235546f[36]),
    .c(al_e6043332),
    .o(al_c665bb87[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ff34e20c (
    .a(ddr_app_wdf_data[37]),
    .b(al_8235546f[37]),
    .c(al_e6043332),
    .o(al_c665bb87[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_16b896f1 (
    .a(ddr_app_wdf_data[38]),
    .b(al_8235546f[38]),
    .c(al_e6043332),
    .o(al_c665bb87[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_6b8db789 (
    .a(ddr_app_wdf_data[39]),
    .b(al_8235546f[39]),
    .c(al_e6043332),
    .o(al_c665bb87[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_39ec6ed3 (
    .a(ddr_app_wdf_data[3]),
    .b(al_8235546f[3]),
    .c(al_e6043332),
    .o(al_c665bb87[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_35940eeb (
    .a(ddr_app_wdf_data[40]),
    .b(al_8235546f[40]),
    .c(al_e6043332),
    .o(al_c665bb87[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b3c61b6c (
    .a(ddr_app_wdf_data[41]),
    .b(al_8235546f[41]),
    .c(al_e6043332),
    .o(al_c665bb87[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_39ff24fb (
    .a(ddr_app_wdf_data[42]),
    .b(al_8235546f[42]),
    .c(al_e6043332),
    .o(al_c665bb87[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9ad6e184 (
    .a(ddr_app_wdf_data[43]),
    .b(al_8235546f[43]),
    .c(al_e6043332),
    .o(al_c665bb87[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3e6b6094 (
    .a(ddr_app_wdf_data[44]),
    .b(al_8235546f[44]),
    .c(al_e6043332),
    .o(al_c665bb87[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3005da87 (
    .a(ddr_app_wdf_data[45]),
    .b(al_8235546f[45]),
    .c(al_e6043332),
    .o(al_c665bb87[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_af12a03a (
    .a(ddr_app_wdf_data[46]),
    .b(al_8235546f[46]),
    .c(al_e6043332),
    .o(al_c665bb87[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e90aaace (
    .a(ddr_app_wdf_data[47]),
    .b(al_8235546f[47]),
    .c(al_e6043332),
    .o(al_c665bb87[47]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5b070695 (
    .a(ddr_app_wdf_data[48]),
    .b(al_8235546f[48]),
    .c(al_e6043332),
    .o(al_c665bb87[48]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7458d34d (
    .a(ddr_app_wdf_data[49]),
    .b(al_8235546f[49]),
    .c(al_e6043332),
    .o(al_c665bb87[49]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c018a428 (
    .a(ddr_app_wdf_data[4]),
    .b(al_8235546f[4]),
    .c(al_e6043332),
    .o(al_c665bb87[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9817f99f (
    .a(ddr_app_wdf_data[50]),
    .b(al_8235546f[50]),
    .c(al_e6043332),
    .o(al_c665bb87[50]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_613ddd7 (
    .a(ddr_app_wdf_data[51]),
    .b(al_8235546f[51]),
    .c(al_e6043332),
    .o(al_c665bb87[51]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_981b85d9 (
    .a(ddr_app_wdf_data[52]),
    .b(al_8235546f[52]),
    .c(al_e6043332),
    .o(al_c665bb87[52]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c9da3e04 (
    .a(ddr_app_wdf_data[53]),
    .b(al_8235546f[53]),
    .c(al_e6043332),
    .o(al_c665bb87[53]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3344f2be (
    .a(ddr_app_wdf_data[54]),
    .b(al_8235546f[54]),
    .c(al_e6043332),
    .o(al_c665bb87[54]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fa72e426 (
    .a(ddr_app_wdf_data[55]),
    .b(al_8235546f[55]),
    .c(al_e6043332),
    .o(al_c665bb87[55]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a15dd36d (
    .a(ddr_app_wdf_data[56]),
    .b(al_8235546f[56]),
    .c(al_e6043332),
    .o(al_c665bb87[56]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2132087b (
    .a(ddr_app_wdf_data[57]),
    .b(al_8235546f[57]),
    .c(al_e6043332),
    .o(al_c665bb87[57]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d3c2f008 (
    .a(ddr_app_wdf_data[58]),
    .b(al_8235546f[58]),
    .c(al_e6043332),
    .o(al_c665bb87[58]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a6ddcc63 (
    .a(ddr_app_wdf_data[59]),
    .b(al_8235546f[59]),
    .c(al_e6043332),
    .o(al_c665bb87[59]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_cbc6406f (
    .a(ddr_app_wdf_data[5]),
    .b(al_8235546f[5]),
    .c(al_e6043332),
    .o(al_c665bb87[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2ca61c64 (
    .a(ddr_app_wdf_data[60]),
    .b(al_8235546f[60]),
    .c(al_e6043332),
    .o(al_c665bb87[60]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_37f72ca2 (
    .a(ddr_app_wdf_data[61]),
    .b(al_8235546f[61]),
    .c(al_e6043332),
    .o(al_c665bb87[61]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5161eab (
    .a(ddr_app_wdf_data[62]),
    .b(al_8235546f[62]),
    .c(al_e6043332),
    .o(al_c665bb87[62]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_25c5c8ad (
    .a(ddr_app_wdf_data[63]),
    .b(al_8235546f[63]),
    .c(al_e6043332),
    .o(al_c665bb87[63]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c8cd9ada (
    .a(ddr_app_wdf_data[64]),
    .b(al_8235546f[64]),
    .c(al_e6043332),
    .o(al_c665bb87[64]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d3e08631 (
    .a(ddr_app_wdf_data[65]),
    .b(al_8235546f[65]),
    .c(al_e6043332),
    .o(al_c665bb87[65]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_6bb9ce25 (
    .a(ddr_app_wdf_data[66]),
    .b(al_8235546f[66]),
    .c(al_e6043332),
    .o(al_c665bb87[66]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7555e3fb (
    .a(ddr_app_wdf_data[67]),
    .b(al_8235546f[67]),
    .c(al_e6043332),
    .o(al_c665bb87[67]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5eae484f (
    .a(ddr_app_wdf_data[68]),
    .b(al_8235546f[68]),
    .c(al_e6043332),
    .o(al_c665bb87[68]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a7f85bd1 (
    .a(ddr_app_wdf_data[69]),
    .b(al_8235546f[69]),
    .c(al_e6043332),
    .o(al_c665bb87[69]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_181f84ca (
    .a(ddr_app_wdf_data[6]),
    .b(al_8235546f[6]),
    .c(al_e6043332),
    .o(al_c665bb87[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_24335f6d (
    .a(ddr_app_wdf_data[70]),
    .b(al_8235546f[70]),
    .c(al_e6043332),
    .o(al_c665bb87[70]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b8d43574 (
    .a(ddr_app_wdf_data[71]),
    .b(al_8235546f[71]),
    .c(al_e6043332),
    .o(al_c665bb87[71]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_823a0576 (
    .a(ddr_app_wdf_data[72]),
    .b(al_8235546f[72]),
    .c(al_e6043332),
    .o(al_c665bb87[72]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_156a082e (
    .a(ddr_app_wdf_data[73]),
    .b(al_8235546f[73]),
    .c(al_e6043332),
    .o(al_c665bb87[73]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2479f4f7 (
    .a(ddr_app_wdf_data[74]),
    .b(al_8235546f[74]),
    .c(al_e6043332),
    .o(al_c665bb87[74]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4912e320 (
    .a(ddr_app_wdf_data[75]),
    .b(al_8235546f[75]),
    .c(al_e6043332),
    .o(al_c665bb87[75]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5e90552b (
    .a(ddr_app_wdf_data[76]),
    .b(al_8235546f[76]),
    .c(al_e6043332),
    .o(al_c665bb87[76]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5f0aab7e (
    .a(ddr_app_wdf_data[77]),
    .b(al_8235546f[77]),
    .c(al_e6043332),
    .o(al_c665bb87[77]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_bc157ba5 (
    .a(ddr_app_wdf_data[78]),
    .b(al_8235546f[78]),
    .c(al_e6043332),
    .o(al_c665bb87[78]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_701ae803 (
    .a(ddr_app_wdf_data[79]),
    .b(al_8235546f[79]),
    .c(al_e6043332),
    .o(al_c665bb87[79]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_75799494 (
    .a(ddr_app_wdf_data[7]),
    .b(al_8235546f[7]),
    .c(al_e6043332),
    .o(al_c665bb87[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f9ce42b3 (
    .a(ddr_app_wdf_data[80]),
    .b(al_8235546f[80]),
    .c(al_e6043332),
    .o(al_c665bb87[80]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3e7a4af6 (
    .a(ddr_app_wdf_data[81]),
    .b(al_8235546f[81]),
    .c(al_e6043332),
    .o(al_c665bb87[81]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_913ecced (
    .a(ddr_app_wdf_data[82]),
    .b(al_8235546f[82]),
    .c(al_e6043332),
    .o(al_c665bb87[82]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ebab35b0 (
    .a(ddr_app_wdf_data[83]),
    .b(al_8235546f[83]),
    .c(al_e6043332),
    .o(al_c665bb87[83]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a5a40575 (
    .a(ddr_app_wdf_data[84]),
    .b(al_8235546f[84]),
    .c(al_e6043332),
    .o(al_c665bb87[84]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7a6b9893 (
    .a(ddr_app_wdf_data[85]),
    .b(al_8235546f[85]),
    .c(al_e6043332),
    .o(al_c665bb87[85]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d687e0fd (
    .a(ddr_app_wdf_data[86]),
    .b(al_8235546f[86]),
    .c(al_e6043332),
    .o(al_c665bb87[86]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7600856e (
    .a(ddr_app_wdf_data[87]),
    .b(al_8235546f[87]),
    .c(al_e6043332),
    .o(al_c665bb87[87]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1ff0bee1 (
    .a(ddr_app_wdf_data[88]),
    .b(al_8235546f[88]),
    .c(al_e6043332),
    .o(al_c665bb87[88]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_205c8e0a (
    .a(ddr_app_wdf_data[89]),
    .b(al_8235546f[89]),
    .c(al_e6043332),
    .o(al_c665bb87[89]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d36db104 (
    .a(ddr_app_wdf_data[8]),
    .b(al_8235546f[8]),
    .c(al_e6043332),
    .o(al_c665bb87[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7043fc55 (
    .a(ddr_app_wdf_data[90]),
    .b(al_8235546f[90]),
    .c(al_e6043332),
    .o(al_c665bb87[90]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b53cc7c5 (
    .a(ddr_app_wdf_data[91]),
    .b(al_8235546f[91]),
    .c(al_e6043332),
    .o(al_c665bb87[91]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e24d3f13 (
    .a(ddr_app_wdf_data[92]),
    .b(al_8235546f[92]),
    .c(al_e6043332),
    .o(al_c665bb87[92]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b78d88f0 (
    .a(ddr_app_wdf_data[93]),
    .b(al_8235546f[93]),
    .c(al_e6043332),
    .o(al_c665bb87[93]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_26022094 (
    .a(ddr_app_wdf_data[94]),
    .b(al_8235546f[94]),
    .c(al_e6043332),
    .o(al_c665bb87[94]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d948091e (
    .a(ddr_app_wdf_data[95]),
    .b(al_8235546f[95]),
    .c(al_e6043332),
    .o(al_c665bb87[95]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c18c5d45 (
    .a(ddr_app_wdf_data[96]),
    .b(al_8235546f[96]),
    .c(al_e6043332),
    .o(al_c665bb87[96]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_29788b90 (
    .a(ddr_app_wdf_data[97]),
    .b(al_8235546f[97]),
    .c(al_e6043332),
    .o(al_c665bb87[97]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d388bf90 (
    .a(ddr_app_wdf_data[98]),
    .b(al_8235546f[98]),
    .c(al_e6043332),
    .o(al_c665bb87[98]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_33e38df4 (
    .a(ddr_app_wdf_data[99]),
    .b(al_8235546f[99]),
    .c(al_e6043332),
    .o(al_c665bb87[99]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9422cc07 (
    .a(ddr_app_wdf_data[9]),
    .b(al_8235546f[9]),
    .c(al_e6043332),
    .o(al_c665bb87[9]));
  AL_DFF_0 al_8b629200 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e837a56c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b7d1c4));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT(16'h2230))
    al_c3449d63 (
    .a(ddr_app_wdf_end),
    .b(al_6db5b9d2),
    .c(al_6b7d1c4),
    .d(al_d872bb7e),
    .o(al_e837a56c));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_27ea7b1e (
    .a(ddr_app_wdf_mask[0]),
    .b(al_eb430c3c[0]),
    .c(al_fd258f8),
    .o(al_e8087d79[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_bf06af26 (
    .a(ddr_app_wdf_mask[10]),
    .b(al_eb430c3c[10]),
    .c(al_fd258f8),
    .o(al_e8087d79[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d5534096 (
    .a(ddr_app_wdf_mask[11]),
    .b(al_eb430c3c[11]),
    .c(al_fd258f8),
    .o(al_e8087d79[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1171172d (
    .a(ddr_app_wdf_mask[12]),
    .b(al_eb430c3c[12]),
    .c(al_fd258f8),
    .o(al_e8087d79[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c0fa9e7 (
    .a(ddr_app_wdf_mask[13]),
    .b(al_eb430c3c[13]),
    .c(al_fd258f8),
    .o(al_e8087d79[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a67a1359 (
    .a(ddr_app_wdf_mask[14]),
    .b(al_eb430c3c[14]),
    .c(al_fd258f8),
    .o(al_e8087d79[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c8e4f6e8 (
    .a(ddr_app_wdf_mask[15]),
    .b(al_eb430c3c[15]),
    .c(al_fd258f8),
    .o(al_e8087d79[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_26964dde (
    .a(ddr_app_wdf_mask[16]),
    .b(al_eb430c3c[16]),
    .c(al_fd258f8),
    .o(al_e8087d79[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9eef0c34 (
    .a(ddr_app_wdf_mask[17]),
    .b(al_eb430c3c[17]),
    .c(al_fd258f8),
    .o(al_e8087d79[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5a0394cf (
    .a(ddr_app_wdf_mask[18]),
    .b(al_eb430c3c[18]),
    .c(al_fd258f8),
    .o(al_e8087d79[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a96f986 (
    .a(ddr_app_wdf_mask[19]),
    .b(al_eb430c3c[19]),
    .c(al_fd258f8),
    .o(al_e8087d79[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_390ace36 (
    .a(ddr_app_wdf_mask[1]),
    .b(al_eb430c3c[1]),
    .c(al_fd258f8),
    .o(al_e8087d79[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_29bda364 (
    .a(ddr_app_wdf_mask[20]),
    .b(al_eb430c3c[20]),
    .c(al_fd258f8),
    .o(al_e8087d79[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1a3f5a76 (
    .a(ddr_app_wdf_mask[21]),
    .b(al_eb430c3c[21]),
    .c(al_fd258f8),
    .o(al_e8087d79[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fc88a5a (
    .a(ddr_app_wdf_mask[22]),
    .b(al_eb430c3c[22]),
    .c(al_fd258f8),
    .o(al_e8087d79[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_496ef5ff (
    .a(ddr_app_wdf_mask[23]),
    .b(al_eb430c3c[23]),
    .c(al_fd258f8),
    .o(al_e8087d79[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_668aed3a (
    .a(ddr_app_wdf_mask[24]),
    .b(al_eb430c3c[24]),
    .c(al_fd258f8),
    .o(al_e8087d79[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1feb3d2e (
    .a(ddr_app_wdf_mask[25]),
    .b(al_eb430c3c[25]),
    .c(al_fd258f8),
    .o(al_e8087d79[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_bebdfe5b (
    .a(ddr_app_wdf_mask[26]),
    .b(al_eb430c3c[26]),
    .c(al_fd258f8),
    .o(al_e8087d79[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4659a630 (
    .a(ddr_app_wdf_mask[27]),
    .b(al_eb430c3c[27]),
    .c(al_fd258f8),
    .o(al_e8087d79[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_6920d2f7 (
    .a(ddr_app_wdf_mask[28]),
    .b(al_eb430c3c[28]),
    .c(al_fd258f8),
    .o(al_e8087d79[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4696ddb9 (
    .a(ddr_app_wdf_mask[29]),
    .b(al_eb430c3c[29]),
    .c(al_fd258f8),
    .o(al_e8087d79[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5ad1f9df (
    .a(ddr_app_wdf_mask[2]),
    .b(al_eb430c3c[2]),
    .c(al_fd258f8),
    .o(al_e8087d79[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_99d8fa03 (
    .a(ddr_app_wdf_mask[30]),
    .b(al_eb430c3c[30]),
    .c(al_fd258f8),
    .o(al_e8087d79[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e7a279e (
    .a(ddr_app_wdf_mask[31]),
    .b(al_eb430c3c[31]),
    .c(al_fd258f8),
    .o(al_e8087d79[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_96d0ee15 (
    .a(ddr_app_wdf_mask[3]),
    .b(al_eb430c3c[3]),
    .c(al_fd258f8),
    .o(al_e8087d79[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ce045dc2 (
    .a(ddr_app_wdf_mask[4]),
    .b(al_eb430c3c[4]),
    .c(al_fd258f8),
    .o(al_e8087d79[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e21787ad (
    .a(ddr_app_wdf_mask[5]),
    .b(al_eb430c3c[5]),
    .c(al_fd258f8),
    .o(al_e8087d79[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_14643808 (
    .a(ddr_app_wdf_mask[6]),
    .b(al_eb430c3c[6]),
    .c(al_fd258f8),
    .o(al_e8087d79[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_bd077f07 (
    .a(ddr_app_wdf_mask[7]),
    .b(al_eb430c3c[7]),
    .c(al_fd258f8),
    .o(al_e8087d79[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8501c24b (
    .a(ddr_app_wdf_mask[8]),
    .b(al_eb430c3c[8]),
    .c(al_fd258f8),
    .o(al_e8087d79[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_3c169a08 (
    .a(ddr_app_wdf_mask[9]),
    .b(al_eb430c3c[9]),
    .c(al_fd258f8),
    .o(al_e8087d79[9]));
  AL_DFF_0 al_78c7dbfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cf2346e1),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_6ab6f142));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_bde808a3 (
    .i(al_6ab6f142),
    .o(al_3daf893a));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9fd64251 (
    .i(al_3daf893a),
    .o(al_947c0ab9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_9b86d42b (
    .i(al_6ab6f142),
    .o(al_2b896d2b));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_44a6811e (
    .i(al_2b896d2b),
    .o(al_e6043332));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1d080d18 (
    .i(al_6ab6f142),
    .o(al_6d2ef296));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7e2afd20 (
    .i(al_6d2ef296),
    .o(al_9431cde9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1537f143 (
    .i(al_6ab6f142),
    .o(al_4fdebbe9));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e6f6ec90 (
    .i(al_4fdebbe9),
    .o(al_b456bf15));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_94c74413 (
    .i(al_6ab6f142),
    .o(al_d56bc9f8));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_591afd5d (
    .i(al_d56bc9f8),
    .o(al_fd258f8));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_accb03d5 (
    .i(al_6ab6f142),
    .o(al_630d6511));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c2998070 (
    .i(al_630d6511),
    .o(al_1ceb77fa));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7a776a42 (
    .i(al_6ab6f142),
    .o(al_ba561a9e));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2c3edb81 (
    .i(al_ba561a9e),
    .o(al_d872bb7e));
  AL_DFF_0 al_178842fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_3021b8d9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5ed629c8));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT(16'h2230))
    al_49596466 (
    .a(ddr_app_wdf_wren),
    .b(al_6db5b9d2),
    .c(al_5ed629c8),
    .d(al_1ceb77fa),
    .o(al_3021b8d9));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_cdce2e8 (
    .a(al_603c814),
    .b(al_2ca0cac1),
    .o(al_2d1611fb));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5561a0da (
    .a(al_af133298[5]),
    .b(al_162fb89b[0]),
    .c(al_f49dc4e0),
    .o(al_1e58d748[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_90006a7e (
    .a(al_af133298[6]),
    .b(al_162fb89b[1]),
    .c(al_f49dc4e0),
    .o(al_1e58d748[1]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_b6bd62b1 (
    .a(al_cc4d831c[1]),
    .b(al_60b9b0f8),
    .o(al_17f22329));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9004739 (
    .di(al_1e58d748),
    .raddr({1'b0,al_cdc129c7}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({1'b0,al_4e964d68[3:0]}),
    .wclk(al_ef3696df[0]),
    .we(al_17f22329),
    .rdo(al_75c0d27f[1:0]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2607ea08 (
    .di(al_1e58d748),
    .raddr({1'b0,al_c394d21b}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({1'b0,al_4e964d68[3:0]}),
    .wclk(al_ef3696df[0]),
    .we(al_17f22329),
    .rdo(al_a2dfc1ad[1:0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8859416b (
    .a(al_af133298[7]),
    .b(al_162fb89b[2]),
    .c(al_f49dc4e0),
    .o(al_98ae77f2[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a33bdf4f (
    .a(al_af133298[8]),
    .b(al_162fb89b[3]),
    .c(al_f49dc4e0),
    .o(al_98ae77f2[1]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_a421f798 (
    .di(al_98ae77f2),
    .raddr({1'b0,al_cdc129c7}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({1'b0,al_4e964d68[3:0]}),
    .wclk(al_ef3696df[0]),
    .we(al_17f22329),
    .rdo(al_75c0d27f[3:2]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_df535c67 (
    .di(al_98ae77f2),
    .raddr({1'b0,al_c394d21b}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({1'b0,al_4e964d68[3:0]}),
    .wclk(al_ef3696df[0]),
    .we(al_17f22329),
    .rdo(al_a2dfc1ad[3:2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_ade67499 (
    .a(al_162fb89b[0]),
    .b(al_f49dc4e0),
    .c(al_57c38d66[0]),
    .o(al_4e964d68[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_443c0b7f (
    .a(al_162fb89b[1]),
    .b(al_f49dc4e0),
    .c(al_57c38d66[1]),
    .o(al_4e964d68[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_59c538f0 (
    .a(al_162fb89b[2]),
    .b(al_f49dc4e0),
    .c(al_57c38d66[2]),
    .o(al_4e964d68[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_8d07d803 (
    .a(al_162fb89b[3]),
    .b(al_f49dc4e0),
    .c(al_57c38d66[3]),
    .o(al_4e964d68[3]));
  AL_DFF_0 al_ca7af301 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_cc4d831c[1]),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_b9b87e33));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_95c38e28 (
    .i(al_b9b87e33),
    .o(al_64b5f594));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d5c87aeb (
    .i(al_64b5f594),
    .o(al_3730b5bd));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_eb2e732b (
    .i(al_b9b87e33),
    .o(al_e4f5976f));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_ff0d3a53 (
    .i(al_e4f5976f),
    .o(al_2ca0cac1));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    al_132b0bd5 (
    .a(al_603c814),
    .b(al_7cd9f06[1]),
    .c(al_2ca0cac1),
    .o(al_a36f4fe4));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_39bf72c (
    .a(al_603c814),
    .b(al_7cd9f06[4]),
    .c(al_7cd9f06[6]),
    .d(al_2ca0cac1),
    .o(al_9056b393));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_938e654d (
    .a(al_603c814),
    .b(al_7cd9f06[6]),
    .c(al_7cd9f06[8]),
    .d(al_2ca0cac1),
    .o(al_a33220fb));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_1b3168ba (
    .a(al_603c814),
    .b(al_7cd9f06[10]),
    .c(al_7cd9f06[12]),
    .d(al_2ca0cac1),
    .o(al_5e51060a));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_38b23e74 (
    .a(al_603c814),
    .b(al_7cd9f06[0]),
    .c(al_7cd9f06[2]),
    .d(al_2ca0cac1),
    .o(al_e0470675));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_6dbfb9f (
    .a(al_603c814),
    .b(al_7cd9f06[5]),
    .c(al_7cd9f06[7]),
    .d(al_2ca0cac1),
    .o(al_44ed9c4));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_2aa28fa5 (
    .a(al_603c814),
    .b(al_7cd9f06[13]),
    .c(al_7cd9f06[15]),
    .d(al_2ca0cac1),
    .o(al_9a26ce4f));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_4714f390 (
    .a(al_603c814),
    .b(al_7cd9f06[1]),
    .c(al_7cd9f06[3]),
    .d(al_2ca0cac1),
    .o(al_1c2bc502));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_532f512f (
    .a(al_603c814),
    .b(al_7cd9f06[11]),
    .c(al_7cd9f06[13]),
    .d(al_2ca0cac1),
    .o(al_aa3cad87));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_bf867686 (
    .a(al_603c814),
    .b(al_7cd9f06[12]),
    .c(al_7cd9f06[14]),
    .d(al_2ca0cac1),
    .o(al_33ae520));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_99c7ca4d (
    .a(al_603c814),
    .b(al_7cd9f06[2]),
    .c(al_7cd9f06[4]),
    .d(al_2ca0cac1),
    .o(al_fba0e4a3));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_4eb7a5f6 (
    .a(al_603c814),
    .b(al_7cd9f06[9]),
    .c(al_7cd9f06[11]),
    .d(al_2ca0cac1),
    .o(al_1fc0eb8a));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_5a32c8b4 (
    .a(al_603c814),
    .b(al_7cd9f06[3]),
    .c(al_7cd9f06[5]),
    .d(al_2ca0cac1),
    .o(al_8a002c3c));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_a2b815cc (
    .a(al_603c814),
    .b(al_7cd9f06[8]),
    .c(al_7cd9f06[10]),
    .d(al_2ca0cac1),
    .o(al_55e87168));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    al_205d13ac (
    .a(al_603c814),
    .b(al_7cd9f06[7]),
    .c(al_7cd9f06[9]),
    .d(al_2ca0cac1),
    .o(al_78b4c22e));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'ha0d8))
    al_f2f4a8a4 (
    .a(al_603c814),
    .b(al_7cd9f06[14]),
    .c(al_7cd9f06[15]),
    .d(al_2ca0cac1),
    .o(al_b8363901));
  AL_DFF_0 al_20cd64d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[0]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[0]));
  AL_DFF_0 al_418aa56a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[1]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[1]));
  AL_DFF_0 al_21b1591d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[2]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[2]));
  AL_DFF_0 al_fb815e3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[3]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[3]));
  AL_DFF_0 al_e29b410d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[4]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[4]));
  AL_DFF_0 al_bb751bbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[5]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[5]));
  AL_DFF_0 al_f96031ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[6]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[6]));
  AL_DFF_0 al_7a21d01f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[7]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[7]));
  AL_DFF_0 al_aada2d43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[8]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[8]));
  AL_DFF_0 al_bbe8618e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[9]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[9]));
  AL_DFF_0 al_6d5ac2f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[10]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[10]));
  AL_DFF_0 al_d2c714b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[11]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[11]));
  AL_DFF_0 al_8bd3a39d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[12]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[12]));
  AL_DFF_0 al_db290250 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[13]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[13]));
  AL_DFF_0 al_a3235130 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[14]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[14]));
  AL_DFF_0 al_19347336 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[15]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[15]));
  AL_DFF_0 al_987b769b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[16]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[16]));
  AL_DFF_0 al_740b0acc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[17]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[17]));
  AL_DFF_0 al_66484b46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[18]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[18]));
  AL_DFF_0 al_1ac53769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[19]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[19]));
  AL_DFF_0 al_dbe82378 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[20]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[20]));
  AL_DFF_0 al_9df4a79c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[21]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[21]));
  AL_DFF_0 al_a89b6c87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[22]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[22]));
  AL_DFF_0 al_4b53df31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[23]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[23]));
  AL_DFF_0 al_5164754f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[24]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[24]));
  AL_DFF_0 al_fc9e5760 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[25]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[25]));
  AL_DFF_0 al_c372100 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[26]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[26]));
  AL_DFF_0 al_adce6dfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[27]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[27]));
  AL_DFF_0 al_1dbe54bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[28]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[28]));
  AL_DFF_0 al_4d51196e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[29]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[29]));
  AL_DFF_0 al_eb2d7740 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[30]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[30]));
  AL_DFF_0 al_11febd05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[31]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[31]));
  AL_DFF_0 al_1bdbc3fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[32]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[32]));
  AL_DFF_0 al_be1d07b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[33]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[33]));
  AL_DFF_0 al_4729f79b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[34]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[34]));
  AL_DFF_0 al_d86a53ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[35]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[35]));
  AL_DFF_0 al_7cbeb266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[36]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[36]));
  AL_DFF_0 al_d4ef3579 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[37]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[37]));
  AL_DFF_0 al_f89ad4b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[38]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[38]));
  AL_DFF_0 al_ef304668 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[39]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[39]));
  AL_DFF_0 al_fdc7425b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[40]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[40]));
  AL_DFF_0 al_8a438395 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[41]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[41]));
  AL_DFF_0 al_3cbfd112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[42]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[42]));
  AL_DFF_0 al_b4cd9df0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[43]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[43]));
  AL_DFF_0 al_54c0a5e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[44]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[44]));
  AL_DFF_0 al_b9560613 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[45]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[45]));
  AL_DFF_0 al_f4e576d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[46]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[46]));
  AL_DFF_0 al_aa625ff4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[47]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[47]));
  AL_DFF_0 al_ff735321 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[48]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[48]));
  AL_DFF_0 al_2d70391a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[49]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[49]));
  AL_DFF_0 al_849d4c8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[50]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[50]));
  AL_DFF_0 al_d9826c37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[51]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[51]));
  AL_DFF_0 al_26f785e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[52]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[52]));
  AL_DFF_0 al_9b14671e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[53]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[53]));
  AL_DFF_0 al_908eb1be (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[54]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[54]));
  AL_DFF_0 al_5a3edcf9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[55]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[55]));
  AL_DFF_0 al_34f39324 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[56]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[56]));
  AL_DFF_0 al_93d5175 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[57]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[57]));
  AL_DFF_0 al_9bfa5930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[58]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[58]));
  AL_DFF_0 al_e130202b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[59]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[59]));
  AL_DFF_0 al_f039053 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[60]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[60]));
  AL_DFF_0 al_b9db6b66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[61]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[61]));
  AL_DFF_0 al_5d747db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[62]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[62]));
  AL_DFF_0 al_ddcb373d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[63]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[63]));
  AL_DFF_0 al_c0abc426 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[64]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[64]));
  AL_DFF_0 al_64f0227d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[65]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[65]));
  AL_DFF_0 al_1f304677 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[66]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[66]));
  AL_DFF_0 al_f9cb2d5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[67]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[67]));
  AL_DFF_0 al_5c0647b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[68]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[68]));
  AL_DFF_0 al_56a62246 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[69]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[69]));
  AL_DFF_0 al_da7555d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[70]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[70]));
  AL_DFF_0 al_34dd34a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[71]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[71]));
  AL_DFF_0 al_fe0ad443 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[72]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[72]));
  AL_DFF_0 al_f94f8435 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[73]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[73]));
  AL_DFF_0 al_ec370534 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[74]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[74]));
  AL_DFF_0 al_21bf312 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[75]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[75]));
  AL_DFF_0 al_fcf161aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[76]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[76]));
  AL_DFF_0 al_f7e89c88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[77]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[77]));
  AL_DFF_0 al_dc5e845a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[78]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[78]));
  AL_DFF_0 al_7b0f188d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[79]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[79]));
  AL_DFF_0 al_fdb3c9eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[80]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[80]));
  AL_DFF_0 al_a009f392 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[81]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[81]));
  AL_DFF_0 al_481362de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[82]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[82]));
  AL_DFF_0 al_5f14e22d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[83]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[83]));
  AL_DFF_0 al_c15ae1cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[84]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[84]));
  AL_DFF_0 al_20a7b873 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[85]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[85]));
  AL_DFF_0 al_ac959197 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[86]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[86]));
  AL_DFF_0 al_9c5aaa0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[87]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[87]));
  AL_DFF_0 al_dda37f2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[88]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[88]));
  AL_DFF_0 al_b64ac06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[89]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[89]));
  AL_DFF_0 al_a33172ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[90]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[90]));
  AL_DFF_0 al_6276107e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[91]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[91]));
  AL_DFF_0 al_28b77b62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[92]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[92]));
  AL_DFF_0 al_a3b1834 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[93]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[93]));
  AL_DFF_0 al_28fcf581 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[94]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[94]));
  AL_DFF_0 al_41c35b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[95]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[95]));
  AL_DFF_0 al_7c97c115 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[96]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[96]));
  AL_DFF_0 al_3d877221 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[97]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[97]));
  AL_DFF_0 al_5e54ba56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[98]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[98]));
  AL_DFF_0 al_2cc71769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[99]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[99]));
  AL_DFF_0 al_782fd1f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[100]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[100]));
  AL_DFF_0 al_a91b680 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[101]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[101]));
  AL_DFF_0 al_745cec3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[102]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[102]));
  AL_DFF_0 al_f7248a09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[103]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[103]));
  AL_DFF_0 al_f1d04629 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[104]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[104]));
  AL_DFF_0 al_c94ac04d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[105]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[105]));
  AL_DFF_0 al_577ba96c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[106]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[106]));
  AL_DFF_0 al_683391de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[107]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[107]));
  AL_DFF_0 al_a410584f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[108]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[108]));
  AL_DFF_0 al_d0cd60b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[109]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[109]));
  AL_DFF_0 al_ecce7582 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[110]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[110]));
  AL_DFF_0 al_edf548a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[111]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[111]));
  AL_DFF_0 al_f913c675 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[112]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[112]));
  AL_DFF_0 al_29dce1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[113]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[113]));
  AL_DFF_0 al_6ec8198c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[114]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[114]));
  AL_DFF_0 al_10b84044 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[115]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[115]));
  AL_DFF_0 al_1f92e8b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[116]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[116]));
  AL_DFF_0 al_3a4377fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[117]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[117]));
  AL_DFF_0 al_e8499953 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[118]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[118]));
  AL_DFF_0 al_fd47d903 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[119]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[119]));
  AL_DFF_0 al_825ffe37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[120]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[120]));
  AL_DFF_0 al_175025fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[121]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[121]));
  AL_DFF_0 al_31a7488 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[122]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[122]));
  AL_DFF_0 al_a33fb79b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[123]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[123]));
  AL_DFF_0 al_e0d33bcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[124]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[124]));
  AL_DFF_0 al_ae200f3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[125]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[125]));
  AL_DFF_0 al_20735b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[126]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[126]));
  AL_DFF_0 al_8bd14c4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[127]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[127]));
  AL_DFF_0 al_db14af65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[128]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[128]));
  AL_DFF_0 al_5fa8ef3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[129]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[129]));
  AL_DFF_0 al_124f8119 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[130]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[130]));
  AL_DFF_0 al_a83c5455 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[131]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[131]));
  AL_DFF_0 al_92bfb0a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[132]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[132]));
  AL_DFF_0 al_74e8bcdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[133]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[133]));
  AL_DFF_0 al_741d36e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[134]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[134]));
  AL_DFF_0 al_1764776c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[135]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[135]));
  AL_DFF_0 al_b35daefe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[136]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[136]));
  AL_DFF_0 al_5fa31781 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[137]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[137]));
  AL_DFF_0 al_11601c9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[138]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[138]));
  AL_DFF_0 al_e3c4cb79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[139]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[139]));
  AL_DFF_0 al_d9539f50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[140]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[140]));
  AL_DFF_0 al_ea5c2b39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[141]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[141]));
  AL_DFF_0 al_49c26606 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[142]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[142]));
  AL_DFF_0 al_c0c79fc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[143]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[143]));
  AL_DFF_0 al_6389f994 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[144]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[144]));
  AL_DFF_0 al_23262d8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[145]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[145]));
  AL_DFF_0 al_d6c87c87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[146]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[146]));
  AL_DFF_0 al_7cefdb4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[147]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[147]));
  AL_DFF_0 al_3600dfd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[148]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[148]));
  AL_DFF_0 al_cf31450b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[149]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[149]));
  AL_DFF_0 al_92c4209f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[150]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[150]));
  AL_DFF_0 al_a7e9e0b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[151]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[151]));
  AL_DFF_0 al_2f7eb575 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[152]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[152]));
  AL_DFF_0 al_bf592181 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[153]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[153]));
  AL_DFF_0 al_751c8a69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[154]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[154]));
  AL_DFF_0 al_a1547557 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[155]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[155]));
  AL_DFF_0 al_52512160 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[156]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[156]));
  AL_DFF_0 al_18ad5478 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[157]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[157]));
  AL_DFF_0 al_4a01f9ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[158]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[158]));
  AL_DFF_0 al_878b121e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[159]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[159]));
  AL_DFF_0 al_ef59f137 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[160]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[160]));
  AL_DFF_0 al_1b3a4faf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[161]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[161]));
  AL_DFF_0 al_bd533d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[162]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[162]));
  AL_DFF_0 al_aa51c307 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[163]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[163]));
  AL_DFF_0 al_435a8464 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[164]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[164]));
  AL_DFF_0 al_ba110179 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[165]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[165]));
  AL_DFF_0 al_9d9d5c59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[166]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[166]));
  AL_DFF_0 al_32c265f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[167]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[167]));
  AL_DFF_0 al_f821e0de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[168]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[168]));
  AL_DFF_0 al_886a0412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[169]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[169]));
  AL_DFF_0 al_6bff20a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[170]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[170]));
  AL_DFF_0 al_28940b34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[171]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[171]));
  AL_DFF_0 al_784de821 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[172]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[172]));
  AL_DFF_0 al_43493f41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[173]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[173]));
  AL_DFF_0 al_7a18e3f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[174]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[174]));
  AL_DFF_0 al_60a2bf4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[175]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[175]));
  AL_DFF_0 al_f17b3de3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[176]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[176]));
  AL_DFF_0 al_118af70a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[177]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[177]));
  AL_DFF_0 al_fb41892e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[178]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[178]));
  AL_DFF_0 al_726be3ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[179]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[179]));
  AL_DFF_0 al_df9a7d3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[180]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[180]));
  AL_DFF_0 al_3d691c5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[181]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[181]));
  AL_DFF_0 al_76c0f858 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[182]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[182]));
  AL_DFF_0 al_388ebca3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[183]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[183]));
  AL_DFF_0 al_3fbc9256 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[184]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[184]));
  AL_DFF_0 al_5f5893fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[185]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[185]));
  AL_DFF_0 al_d454a920 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[186]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[186]));
  AL_DFF_0 al_cff7e89f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[187]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[187]));
  AL_DFF_0 al_a8b23f94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[188]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[188]));
  AL_DFF_0 al_224b848b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[189]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[189]));
  AL_DFF_0 al_7f08f20e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[190]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[190]));
  AL_DFF_0 al_80c178c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[191]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[191]));
  AL_DFF_0 al_9c1ad667 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[192]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[192]));
  AL_DFF_0 al_56059f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[193]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[193]));
  AL_DFF_0 al_b7ec47eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[194]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[194]));
  AL_DFF_0 al_45eeb7e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[195]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[195]));
  AL_DFF_0 al_df01be6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[196]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[196]));
  AL_DFF_0 al_11f26068 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[197]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[197]));
  AL_DFF_0 al_505214bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[198]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[198]));
  AL_DFF_0 al_e4572915 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[199]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[199]));
  AL_DFF_0 al_d373f9fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[200]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[200]));
  AL_DFF_0 al_c5935e2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[201]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[201]));
  AL_DFF_0 al_94eea95e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[202]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[202]));
  AL_DFF_0 al_57072bea (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[203]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[203]));
  AL_DFF_0 al_4d08d6fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[204]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[204]));
  AL_DFF_0 al_b67365b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[205]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[205]));
  AL_DFF_0 al_fe73f4e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[206]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[206]));
  AL_DFF_0 al_ed6df11e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[207]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[207]));
  AL_DFF_0 al_a0793d10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[208]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[208]));
  AL_DFF_0 al_455deee4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[209]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[209]));
  AL_DFF_0 al_bd5993ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[210]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[210]));
  AL_DFF_0 al_47b12c7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[211]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[211]));
  AL_DFF_0 al_14c8c0fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[212]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[212]));
  AL_DFF_0 al_3b61464d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[213]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[213]));
  AL_DFF_0 al_b26cd948 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[214]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[214]));
  AL_DFF_0 al_aff47cdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[215]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[215]));
  AL_DFF_0 al_7fa78792 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[216]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[216]));
  AL_DFF_0 al_42f3ebbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[217]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[217]));
  AL_DFF_0 al_ac23e58d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[218]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[218]));
  AL_DFF_0 al_a6c11b8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[219]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[219]));
  AL_DFF_0 al_38186f85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[220]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[220]));
  AL_DFF_0 al_c3f592a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[221]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[221]));
  AL_DFF_0 al_92dfee6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[222]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[222]));
  AL_DFF_0 al_33bf3e6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[223]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[223]));
  AL_DFF_0 al_14402954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[224]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[224]));
  AL_DFF_0 al_9e76c5fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[225]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[225]));
  AL_DFF_0 al_38bb9081 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[226]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[226]));
  AL_DFF_0 al_ae4a1ffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[227]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[227]));
  AL_DFF_0 al_1033b729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[228]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[228]));
  AL_DFF_0 al_ca4ec8c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[229]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[229]));
  AL_DFF_0 al_24cc8962 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[230]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[230]));
  AL_DFF_0 al_d4b627fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[231]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[231]));
  AL_DFF_0 al_d47bc4ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[232]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[232]));
  AL_DFF_0 al_22281262 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[233]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[233]));
  AL_DFF_0 al_1d092166 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[234]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[234]));
  AL_DFF_0 al_769a277f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[235]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[235]));
  AL_DFF_0 al_92def549 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[236]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[236]));
  AL_DFF_0 al_1d7f490 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[237]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[237]));
  AL_DFF_0 al_ebfd0e6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[238]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[238]));
  AL_DFF_0 al_6691d8c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[239]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[239]));
  AL_DFF_0 al_5d8d5baa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[240]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[240]));
  AL_DFF_0 al_88784f6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[241]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[241]));
  AL_DFF_0 al_c689dcb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[242]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[242]));
  AL_DFF_0 al_20692ea8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[243]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[243]));
  AL_DFF_0 al_4cc15d5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[244]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[244]));
  AL_DFF_0 al_16aeb2d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[245]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[245]));
  AL_DFF_0 al_febf7708 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[246]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[246]));
  AL_DFF_0 al_7b28cca4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[247]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[247]));
  AL_DFF_0 al_10b6561e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[248]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[248]));
  AL_DFF_0 al_e2d540b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[249]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[249]));
  AL_DFF_0 al_9f6a0510 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[250]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[250]));
  AL_DFF_0 al_6a64aca8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[251]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[251]));
  AL_DFF_0 al_47d7303 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[252]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[252]));
  AL_DFF_0 al_cd466662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[253]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[253]));
  AL_DFF_0 al_a8a4cfbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[254]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[254]));
  AL_DFF_0 al_c3a9debc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_data[255]),
    .en(al_e6043332),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8235546f[255]));
  AL_DFF_0 al_db4ee810 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[0]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[0]));
  AL_DFF_0 al_ea3a0e4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[1]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[1]));
  AL_DFF_0 al_ee3131fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[2]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[2]));
  AL_DFF_0 al_f4608d2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[3]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[3]));
  AL_DFF_0 al_bd3fc19f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[4]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[4]));
  AL_DFF_0 al_ef6a5690 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[5]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[5]));
  AL_DFF_0 al_71bbb086 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[6]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[6]));
  AL_DFF_0 al_d422dd72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[7]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[7]));
  AL_DFF_0 al_917e75dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[8]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[8]));
  AL_DFF_0 al_a6c2873f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[9]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[9]));
  AL_DFF_0 al_5e809a9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[10]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[10]));
  AL_DFF_0 al_f7458b99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[11]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[11]));
  AL_DFF_0 al_8e2e5190 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[12]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[12]));
  AL_DFF_0 al_31be4661 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[13]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[13]));
  AL_DFF_0 al_51cabcfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[14]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[14]));
  AL_DFF_0 al_1b5f8112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[15]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[15]));
  AL_DFF_0 al_c0f95ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[16]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[16]));
  AL_DFF_0 al_38d08417 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[17]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[17]));
  AL_DFF_0 al_4bc222a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[18]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[18]));
  AL_DFF_0 al_6af8f126 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[19]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[19]));
  AL_DFF_0 al_873e976a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[20]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[20]));
  AL_DFF_0 al_2cbc584d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[21]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[21]));
  AL_DFF_0 al_d2933792 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[22]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[22]));
  AL_DFF_0 al_8216a9da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[23]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[23]));
  AL_DFF_0 al_fed62540 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[24]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[24]));
  AL_DFF_0 al_3848e910 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[25]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[25]));
  AL_DFF_0 al_21cd416b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[26]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[26]));
  AL_DFF_0 al_cdc61820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[27]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[27]));
  AL_DFF_0 al_619393e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[28]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[28]));
  AL_DFF_0 al_147eb6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[29]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[29]));
  AL_DFF_0 al_5e41258e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[30]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[30]));
  AL_DFF_0 al_1f5bff71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(ddr_app_wdf_mask[31]),
    .en(al_fd258f8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb430c3c[31]));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_aafc25f7 (
    .a(al_1308b999),
    .b(al_6db5b9d2),
    .c(al_cdc129c7[0]),
    .d(al_cdc129c7[1]),
    .e(al_cdc129c7[2]),
    .o(al_f9e997a5));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_f2275f83 (
    .a(al_1308b999),
    .b(al_6db5b9d2),
    .c(al_cdc129c7[0]),
    .d(al_cdc129c7[1]),
    .o(al_f24aaa07));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_74c63ac8 (
    .a(al_1308b999),
    .b(al_6db5b9d2),
    .c(al_cdc129c7[0]),
    .o(al_984d7f7));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_f8b65bd0 (
    .a(al_1308b999),
    .b(al_6db5b9d2),
    .c(al_cdc129c7[0]),
    .d(al_cdc129c7[1]),
    .e(al_cdc129c7[2]),
    .f(al_cdc129c7[3]),
    .o(al_1819221f));
  AL_DFF_0 al_6e21997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_984d7f7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdc129c7[0]));
  AL_DFF_0 al_b4cbca1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f24aaa07),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdc129c7[1]));
  AL_DFF_0 al_eccb5156 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_f9e997a5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdc129c7[2]));
  AL_DFF_0 al_716f3664 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1819221f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdc129c7[3]));
  AL_DFF_0 al_2549c526 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a36f4fe4),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[0]));
  AL_DFF_0 al_bee0c765 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_e0470675),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[1]));
  AL_DFF_0 al_b9ad03dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1c2bc502),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[2]));
  AL_DFF_0 al_f92c3ab2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_fba0e4a3),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[3]));
  AL_DFF_0 al_d0f4e1ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8a002c3c),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[4]));
  AL_DFF_0 al_e8044616 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9056b393),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[5]));
  AL_DFF_0 al_53db8e98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44ed9c4),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[6]));
  AL_DFF_0 al_fc46280a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a33220fb),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[7]));
  AL_DFF_0 al_f6d34fc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_78b4c22e),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[8]));
  AL_DFF_0 al_91f3c293 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_55e87168),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[9]));
  AL_DFF_0 al_d34c4876 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_1fc0eb8a),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[10]));
  AL_DFF_0 al_9f6ff8ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_5e51060a),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[11]));
  AL_DFF_0 al_bbcb2548 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_aa3cad87),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[12]));
  AL_DFF_0 al_b052f806 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_33ae520),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[13]));
  AL_DFF_0 al_fa8342c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_9a26ce4f),
    .en(al_2d1611fb),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[14]));
  AL_DFF_0 al_602656b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_b8363901),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7cd9f06[15]));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_57b9d2bd (
    .a(al_cc4d831c[1]),
    .b(al_6db5b9d2),
    .c(al_57c38d66[0]),
    .o(al_555b330b));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_219913be (
    .a(al_cc4d831c[1]),
    .b(al_6db5b9d2),
    .c(al_57c38d66[0]),
    .d(al_57c38d66[1]),
    .o(al_44a10d10));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_eed0f275 (
    .a(al_cc4d831c[1]),
    .b(al_6db5b9d2),
    .c(al_57c38d66[0]),
    .d(al_57c38d66[1]),
    .e(al_57c38d66[2]),
    .o(al_555cabbf));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_133f0d03 (
    .a(al_cc4d831c[1]),
    .b(al_6db5b9d2),
    .c(al_57c38d66[0]),
    .d(al_57c38d66[1]),
    .e(al_57c38d66[2]),
    .f(al_57c38d66[3]),
    .o(al_8f3c4595));
  AL_DFF_0 al_86453c85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_555b330b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57c38d66[0]));
  AL_DFF_0 al_b99da77c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_44a10d10),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57c38d66[1]));
  AL_DFF_0 al_dc2ab50b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_555cabbf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57c38d66[2]));
  AL_DFF_0 al_d2ab99c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8f3c4595),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57c38d66[3]));
  AL_DFF_0 al_4abf225c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a2dfc1ad[0]),
    .en(al_d22a1e42),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_e0201a[1]));
  AL_DFF_0 al_d01c1ee0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a2dfc1ad[1]),
    .en(al_d22a1e42),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_e0201a[2]));
  AL_DFF_0 al_83d83ba1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a2dfc1ad[2]),
    .en(al_d22a1e42),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_e0201a[3]));
  AL_DFF_0 al_268820db (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a2dfc1ad[3]),
    .en(al_d22a1e42),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_e0201a[4]));
  AL_DFF_0 al_92429166 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[0]));
  AL_DFF_0 al_49d47e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[1]));
  AL_DFF_0 al_2fa70d7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[2]));
  AL_DFF_0 al_a7a504bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[3]));
  AL_DFF_0 al_2caaa353 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[4]));
  AL_DFF_0 al_467dcd6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[5]));
  AL_DFF_0 al_88495593 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[6]));
  AL_DFF_0 al_fab4f51d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[7]));
  AL_DFF_0 al_79494151 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[8]));
  AL_DFF_0 al_c4b1a9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[9]));
  AL_DFF_0 al_80cbd5bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[10]));
  AL_DFF_0 al_a224fc5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[11]));
  AL_DFF_0 al_12298978 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[12]));
  AL_DFF_0 al_97d230d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[13]));
  AL_DFF_0 al_ccf01c9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[14]));
  AL_DFF_0 al_58266b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[15]));
  AL_DFF_0 al_39dd066f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[16]));
  AL_DFF_0 al_2ee6b471 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[17]));
  AL_DFF_0 al_c65ec94a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[18]));
  AL_DFF_0 al_fb9ab0e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[19]));
  AL_DFF_0 al_605061c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[20]));
  AL_DFF_0 al_9b179674 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[21]));
  AL_DFF_0 al_2cc1764e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[22]));
  AL_DFF_0 al_5124461f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[23]));
  AL_DFF_0 al_65284ccf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[24]));
  AL_DFF_0 al_80ca4a72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[25]));
  AL_DFF_0 al_bd1c1acb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[26]));
  AL_DFF_0 al_8cda77d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[27]));
  AL_DFF_0 al_3bab2e85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[28]));
  AL_DFF_0 al_aefa2e89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[29]));
  AL_DFF_0 al_63ef7661 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[30]));
  AL_DFF_0 al_658a4db2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[31]));
  AL_DFF_0 al_c77c49cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[32]));
  AL_DFF_0 al_7736a52c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[33]));
  AL_DFF_0 al_505e4b09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[34]));
  AL_DFF_0 al_7e623c4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[35]));
  AL_DFF_0 al_a54fb72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[36]));
  AL_DFF_0 al_82d5e42e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[37]));
  AL_DFF_0 al_65b56af3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[38]));
  AL_DFF_0 al_8e605d9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[39]));
  AL_DFF_0 al_1fb6e729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[40]));
  AL_DFF_0 al_49c1fecf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[41]));
  AL_DFF_0 al_79948a7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[42]));
  AL_DFF_0 al_3ba99ef2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[43]));
  AL_DFF_0 al_17ca1acb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[44]));
  AL_DFF_0 al_918d11ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[45]));
  AL_DFF_0 al_e2a135c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[46]));
  AL_DFF_0 al_f471dbe6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[47]));
  AL_DFF_0 al_40e13af0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[48]));
  AL_DFF_0 al_34eb21c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[49]));
  AL_DFF_0 al_795a7313 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[50]));
  AL_DFF_0 al_5b1da54a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[51]));
  AL_DFF_0 al_3094e6ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[52]));
  AL_DFF_0 al_406c0ace (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[53]));
  AL_DFF_0 al_fb9fe2f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[54]));
  AL_DFF_0 al_a83678b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[55]));
  AL_DFF_0 al_7b47026b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[56]));
  AL_DFF_0 al_8f33f33f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[57]));
  AL_DFF_0 al_c31097fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[58]));
  AL_DFF_0 al_680cee1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[59]));
  AL_DFF_0 al_39042de9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[60]));
  AL_DFF_0 al_4def353f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[61]));
  AL_DFF_0 al_2fbf159b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[62]));
  AL_DFF_0 al_4287128e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[63]));
  AL_DFF_0 al_748e26d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[64]));
  AL_DFF_0 al_b1aae385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[65]));
  AL_DFF_0 al_e05de010 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[66]));
  AL_DFF_0 al_bfe7efe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[67]));
  AL_DFF_0 al_131459f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[68]));
  AL_DFF_0 al_614c1597 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[69]));
  AL_DFF_0 al_74a5f72c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[70]));
  AL_DFF_0 al_4b240875 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[71]));
  AL_DFF_0 al_131148bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[72]));
  AL_DFF_0 al_68e0ec65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[73]));
  AL_DFF_0 al_8086812f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[74]));
  AL_DFF_0 al_eb66366e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[75]));
  AL_DFF_0 al_a9e25942 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[76]));
  AL_DFF_0 al_4870adbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[77]));
  AL_DFF_0 al_bb8004de (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[78]));
  AL_DFF_0 al_41f05e53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[79]));
  AL_DFF_0 al_bc29a8f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[80]));
  AL_DFF_0 al_94d59b60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[81]));
  AL_DFF_0 al_3547dcf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[82]));
  AL_DFF_0 al_591e42b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[83]));
  AL_DFF_0 al_15523c46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[84]));
  AL_DFF_0 al_efd5b3bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[85]));
  AL_DFF_0 al_2c226eae (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[86]));
  AL_DFF_0 al_4ecda461 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[87]));
  AL_DFF_0 al_b09cf51d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[88]));
  AL_DFF_0 al_67b798c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[89]));
  AL_DFF_0 al_a80c94f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[90]));
  AL_DFF_0 al_173877bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[91]));
  AL_DFF_0 al_f88eabcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[92]));
  AL_DFF_0 al_fd040822 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[93]));
  AL_DFF_0 al_ca90007c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[94]));
  AL_DFF_0 al_de37c937 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[95]));
  AL_DFF_0 al_d4e6f6c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[96]));
  AL_DFF_0 al_3851c62d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[97]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[97]));
  AL_DFF_0 al_f61d44b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[98]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[98]));
  AL_DFF_0 al_1ddcfc2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[99]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[99]));
  AL_DFF_0 al_6d4ac322 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[100]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[100]));
  AL_DFF_0 al_ed28a6c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[101]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[101]));
  AL_DFF_0 al_2262571a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[102]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[102]));
  AL_DFF_0 al_ee4b65b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[103]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[103]));
  AL_DFF_0 al_aa268ff3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[104]));
  AL_DFF_0 al_79bc9092 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[105]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[105]));
  AL_DFF_0 al_92d35f07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[106]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[106]));
  AL_DFF_0 al_a878bed4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[107]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[107]));
  AL_DFF_0 al_95e7c1d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[108]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[108]));
  AL_DFF_0 al_a9454a7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[109]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[109]));
  AL_DFF_0 al_1a90985e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[110]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[110]));
  AL_DFF_0 al_af3a99c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[111]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[111]));
  AL_DFF_0 al_193f361c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[112]));
  AL_DFF_0 al_73ca4c81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[113]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[113]));
  AL_DFF_0 al_6fadaa82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[114]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[114]));
  AL_DFF_0 al_57de020b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[115]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[115]));
  AL_DFF_0 al_e058849d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[116]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[116]));
  AL_DFF_0 al_44de38b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[117]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[117]));
  AL_DFF_0 al_129afb71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[118]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[118]));
  AL_DFF_0 al_21a15bdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[119]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[119]));
  AL_DFF_0 al_d929fca3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[120]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[120]));
  AL_DFF_0 al_172a5753 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[121]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[121]));
  AL_DFF_0 al_dbc2c81a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[122]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[122]));
  AL_DFF_0 al_baba3aac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[123]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[123]));
  AL_DFF_0 al_90fa44d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[124]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[124]));
  AL_DFF_0 al_28632bd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[125]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[125]));
  AL_DFF_0 al_5398a326 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[126]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[126]));
  AL_DFF_0 al_8a89f9e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[127]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[127]));
  AL_DFF_0 al_fb671028 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[128]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[128]));
  AL_DFF_0 al_d037baf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[129]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[129]));
  AL_DFF_0 al_8f7b6057 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[130]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[130]));
  AL_DFF_0 al_5aae87fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[131]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[131]));
  AL_DFF_0 al_e1a7ae70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[132]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[132]));
  AL_DFF_0 al_e18c98f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[133]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[133]));
  AL_DFF_0 al_8c7ca1a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[134]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[134]));
  AL_DFF_0 al_750bbb2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[135]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[135]));
  AL_DFF_0 al_fc6eecdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[136]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[136]));
  AL_DFF_0 al_66f60b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[137]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[137]));
  AL_DFF_0 al_8accff72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[138]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[138]));
  AL_DFF_0 al_4a7f7ec2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[139]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[139]));
  AL_DFF_0 al_e84f4987 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[140]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[140]));
  AL_DFF_0 al_cc817c69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[141]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[141]));
  AL_DFF_0 al_b9c000ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[142]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[142]));
  AL_DFF_0 al_b46ed93b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[143]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[143]));
  AL_DFF_0 al_8e5ec836 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[144]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[144]));
  AL_DFF_0 al_b2f724d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[145]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[145]));
  AL_DFF_0 al_f1c24837 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[146]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[146]));
  AL_DFF_0 al_1941e0ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[147]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[147]));
  AL_DFF_0 al_1d8a7374 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[148]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[148]));
  AL_DFF_0 al_e49365d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[149]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[149]));
  AL_DFF_0 al_744ce86d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[150]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[150]));
  AL_DFF_0 al_16caa2dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[151]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[151]));
  AL_DFF_0 al_9d5c2976 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[152]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[152]));
  AL_DFF_0 al_1375ab46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[153]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[153]));
  AL_DFF_0 al_cbca86be (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[154]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[154]));
  AL_DFF_0 al_61f49746 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[155]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[155]));
  AL_DFF_0 al_42563f92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[156]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[156]));
  AL_DFF_0 al_5affbd58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[157]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[157]));
  AL_DFF_0 al_4f74922b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[158]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[158]));
  AL_DFF_0 al_1993f11d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[159]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[159]));
  AL_DFF_0 al_3a1ffaa3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[160]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[160]));
  AL_DFF_0 al_d6e94857 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[161]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[161]));
  AL_DFF_0 al_3ff1c846 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[162]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[162]));
  AL_DFF_0 al_6817d7f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[163]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[163]));
  AL_DFF_0 al_2dbed35c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[164]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[164]));
  AL_DFF_0 al_b3fbacb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[165]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[165]));
  AL_DFF_0 al_c9a894ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[166]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[166]));
  AL_DFF_0 al_b3e09307 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[167]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[167]));
  AL_DFF_0 al_ba3fcaaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[168]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[168]));
  AL_DFF_0 al_dc8f95e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[169]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[169]));
  AL_DFF_0 al_80b5879d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[170]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[170]));
  AL_DFF_0 al_573b8fa8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[171]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[171]));
  AL_DFF_0 al_f4639d7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[172]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[172]));
  AL_DFF_0 al_edbea8ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[173]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[173]));
  AL_DFF_0 al_ab9f646b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[174]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[174]));
  AL_DFF_0 al_aeeb04b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[175]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[175]));
  AL_DFF_0 al_ddce4a70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[176]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[176]));
  AL_DFF_0 al_37d298fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[177]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[177]));
  AL_DFF_0 al_452ba278 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[178]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[178]));
  AL_DFF_0 al_30e505da (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[179]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[179]));
  AL_DFF_0 al_d9b7c9f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[180]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[180]));
  AL_DFF_0 al_353a7e20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[181]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[181]));
  AL_DFF_0 al_2a38ddf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[182]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[182]));
  AL_DFF_0 al_bdb603b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[183]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[183]));
  AL_DFF_0 al_7e3d5d18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[184]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[184]));
  AL_DFF_0 al_729d526c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[185]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[185]));
  AL_DFF_0 al_6534f94e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[186]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[186]));
  AL_DFF_0 al_e3d94301 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[187]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[187]));
  AL_DFF_0 al_7ef36ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[188]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[188]));
  AL_DFF_0 al_ce98df71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[189]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[189]));
  AL_DFF_0 al_de793dd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[190]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[190]));
  AL_DFF_0 al_599b094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[191]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[191]));
  AL_DFF_0 al_c1397e47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[192]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[192]));
  AL_DFF_0 al_ca4b4025 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[193]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[193]));
  AL_DFF_0 al_6b22f880 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[194]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[194]));
  AL_DFF_0 al_a3965914 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[195]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[195]));
  AL_DFF_0 al_8f6ebe24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[196]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[196]));
  AL_DFF_0 al_6116383f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[197]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[197]));
  AL_DFF_0 al_79ac8c51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[198]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[198]));
  AL_DFF_0 al_8e59f1ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[199]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[199]));
  AL_DFF_0 al_37f5c038 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[200]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[200]));
  AL_DFF_0 al_366bcd35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[201]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[201]));
  AL_DFF_0 al_8a608aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[202]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[202]));
  AL_DFF_0 al_e0c2de3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[203]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[203]));
  AL_DFF_0 al_c784c604 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[204]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[204]));
  AL_DFF_0 al_72e07cf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[205]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[205]));
  AL_DFF_0 al_4254d153 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[206]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[206]));
  AL_DFF_0 al_6f323042 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[207]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[207]));
  AL_DFF_0 al_56dd2e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[208]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[208]));
  AL_DFF_0 al_aef0b80e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[209]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[209]));
  AL_DFF_0 al_908a5c32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[210]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[210]));
  AL_DFF_0 al_a878165c (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[211]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[211]));
  AL_DFF_0 al_86c14cdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[212]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[212]));
  AL_DFF_0 al_5bcf382e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[213]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[213]));
  AL_DFF_0 al_d4ddaff1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[214]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[214]));
  AL_DFF_0 al_627b014f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[215]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[215]));
  AL_DFF_0 al_de724671 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[216]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[216]));
  AL_DFF_0 al_7ed3ba2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[217]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[217]));
  AL_DFF_0 al_2e76cca7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[218]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[218]));
  AL_DFF_0 al_3fd24690 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[219]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[219]));
  AL_DFF_0 al_2c10c04d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[220]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[220]));
  AL_DFF_0 al_4cd0f516 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[221]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[221]));
  AL_DFF_0 al_9a2d1018 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[222]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[222]));
  AL_DFF_0 al_39663de5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[223]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[223]));
  AL_DFF_0 al_1550127f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[224]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[224]));
  AL_DFF_0 al_1bf8e42a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[225]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[225]));
  AL_DFF_0 al_2983e1c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[226]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[226]));
  AL_DFF_0 al_769c661a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[227]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[227]));
  AL_DFF_0 al_b97afa81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[228]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[228]));
  AL_DFF_0 al_4ce8445 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[229]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[229]));
  AL_DFF_0 al_8624f546 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[230]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[230]));
  AL_DFF_0 al_d56d2ab5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[231]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[231]));
  AL_DFF_0 al_8845f480 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[232]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[232]));
  AL_DFF_0 al_27855dff (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[233]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[233]));
  AL_DFF_0 al_2c7626d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[234]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[234]));
  AL_DFF_0 al_dc062730 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[235]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[235]));
  AL_DFF_0 al_abec133 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[236]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[236]));
  AL_DFF_0 al_86f60cc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[237]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[237]));
  AL_DFF_0 al_fc7f298 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[238]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[238]));
  AL_DFF_0 al_df17e2e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[239]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[239]));
  AL_DFF_0 al_56570b54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[240]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[240]));
  AL_DFF_0 al_6068947f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[241]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[241]));
  AL_DFF_0 al_61f1d80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[242]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[242]));
  AL_DFF_0 al_78bcc690 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[243]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[243]));
  AL_DFF_0 al_b9778da1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[244]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[244]));
  AL_DFF_0 al_5f90e4e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[245]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[245]));
  AL_DFF_0 al_b26e1c6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[246]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[246]));
  AL_DFF_0 al_7c5ee836 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[247]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[247]));
  AL_DFF_0 al_2fe9a042 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[248]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[248]));
  AL_DFF_0 al_51fd566e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[249]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[249]));
  AL_DFF_0 al_fc554232 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[250]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[250]));
  AL_DFF_0 al_83d6d835 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[251]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[251]));
  AL_DFF_0 al_2c3e4b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[252]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[252]));
  AL_DFF_0 al_10cc3a1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[253]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[253]));
  AL_DFF_0 al_b535eebf (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[254]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[254]));
  AL_DFF_0 al_2ac58ef3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[255]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[255]));
  AL_DFF_0 al_427027d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[256]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[256]));
  AL_DFF_0 al_8e4e156 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[257]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[257]));
  AL_DFF_0 al_c87335f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[258]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[258]));
  AL_DFF_0 al_1d8e0409 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[259]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[259]));
  AL_DFF_0 al_3a465c84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[260]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[260]));
  AL_DFF_0 al_cf3218ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[261]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[261]));
  AL_DFF_0 al_160e8394 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[262]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[262]));
  AL_DFF_0 al_7ecb461a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[263]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[263]));
  AL_DFF_0 al_6f695116 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[264]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[264]));
  AL_DFF_0 al_f9cc68a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[265]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[265]));
  AL_DFF_0 al_7fa6a79e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[266]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[266]));
  AL_DFF_0 al_81220246 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[267]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[267]));
  AL_DFF_0 al_52e82303 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[268]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[268]));
  AL_DFF_0 al_8600ed00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[269]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[269]));
  AL_DFF_0 al_d20c5ac5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[270]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[270]));
  AL_DFF_0 al_544e78d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[271]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[271]));
  AL_DFF_0 al_984643af (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[272]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[272]));
  AL_DFF_0 al_48193d93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[273]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[273]));
  AL_DFF_0 al_816304e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[274]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[274]));
  AL_DFF_0 al_c2192828 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[275]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[275]));
  AL_DFF_0 al_3cdebf01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[276]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[276]));
  AL_DFF_0 al_eda330b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[277]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[277]));
  AL_DFF_0 al_6101731b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[278]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[278]));
  AL_DFF_0 al_60ea523 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[279]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[279]));
  AL_DFF_0 al_9d8fa271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[280]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[280]));
  AL_DFF_0 al_439e629f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[281]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[281]));
  AL_DFF_0 al_69d27366 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[282]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[282]));
  AL_DFF_0 al_1bf2c51f (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[283]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[283]));
  AL_DFF_0 al_6fe9ff09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[284]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[284]));
  AL_DFF_0 al_1f222d9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[285]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[285]));
  AL_DFF_0 al_406287ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[286]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[286]));
  AL_DFF_0 al_d1820a40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_8c7bed02[287]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e0d53ab[287]));
  AL_DFF_0 al_406492f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f66965[1]),
    .en(al_d22a1e42),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_c394d21b[1]));
  AL_DFF_0 al_5c9c6550 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f66965[2]),
    .en(al_d22a1e42),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_c394d21b[2]));
  AL_DFF_0 al_d5289eb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f66965[3]),
    .en(al_d22a1e42),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_c394d21b[3]));
  AL_DFF_1 al_8656953 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_a3f66965[0]),
    .en(al_d22a1e42),
    .sr(1'b0),
    .ss(al_6db5b9d2),
    .q(al_c394d21b[0]));
  AL_DFF_0 al_17549b69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d1db9874[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3014f961[3]));
  AL_DFF_0 al_56e2777e (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d1db9874[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3014f961[4]));
  AL_DFF_0 al_83b40e3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d1db9874[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3014f961[0]));
  AL_DFF_0 al_764a1e3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d1db9874[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3014f961[1]));
  AL_DFF_0 al_62a0d487 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_d1db9874[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3014f961[2]));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h7430))
    al_12e042b7 (
    .a(al_6b7d1c4),
    .b(al_5ed629c8),
    .c(al_7bc48670),
    .d(al_9431cde9),
    .o(al_6c6fd169));
  AL_DFF_0 al_b0233869 (
    .ar(1'b0),
    .as(1'b0),
    .clk(al_ef3696df[0]),
    .d(al_6c6fd169),
    .en(1'b1),
    .sr(al_6db5b9d2),
    .ss(1'b0),
    .q(al_7bc48670));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    al_8d92153 (
    .a(al_d22a1e42),
    .b(al_6db5b9d2),
    .c(al_e0201a[1]),
    .d(al_a2dfc1ad[0]),
    .o(al_9c7fabce[1]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    al_50219b78 (
    .a(al_d22a1e42),
    .b(al_6db5b9d2),
    .c(al_e0201a[2]),
    .d(al_a2dfc1ad[1]),
    .o(al_9c7fabce[2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    al_27f9ee61 (
    .a(al_d22a1e42),
    .b(al_6db5b9d2),
    .c(al_e0201a[3]),
    .d(al_a2dfc1ad[2]),
    .o(al_9c7fabce[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_edb94000 (
    .a(al_6b7d1c4),
    .b(al_5ed629c8),
    .c(al_947c0ab9),
    .o(al_603c814));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~E*~(~D*~(C*A))))"),
    .INIT(32'hcccc004c))
    al_dbbc376 (
    .a(al_603c814),
    .b(al_eaa97ed5),
    .c(al_7cd9f06[14]),
    .d(al_7cd9f06[15]),
    .e(al_2ca0cac1),
    .o(al_cf2346e1));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~C)*~(B*A))"),
    .INIT(16'h8f88))
    al_597cdf2e (
    .a(al_cf2346e1),
    .b(al_603c814),
    .c(al_b456bf15),
    .d(al_2ca0cac1),
    .o(al_d22a1e42));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    al_c46d42a0 (
    .a(al_d22a1e42),
    .b(al_6db5b9d2),
    .c(al_e0201a[4]),
    .d(al_a2dfc1ad[3]),
    .o(al_9c7fabce[4]));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~E*~(~D*~(C*A))))"),
    .INIT(32'hcccc004c))
    al_1cc0570 (
    .a(al_603c814),
    .b(al_2acf9590),
    .c(al_7cd9f06[14]),
    .d(al_7cd9f06[15]),
    .e(al_3730b5bd),
    .o(al_b03fffe1));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d46df3fd (
    .di(al_c665bb87[5:4]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[5:4]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7e0d19c8 (
    .di(al_c665bb87[3:2]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[3:2]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_eff53562 (
    .di(al_c665bb87[1:0]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[1:0]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_1a312f0e (
    .di(al_c665bb87[65:64]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[65:64]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_8b5a1672 (
    .di(al_c665bb87[63:62]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[63:62]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b9c4f88f (
    .di(al_c665bb87[61:60]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[61:60]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_96b5c388 (
    .di(al_c665bb87[71:70]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[71:70]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2d3b0023 (
    .di(al_c665bb87[69:68]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[69:68]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7ae8df5c (
    .di(al_c665bb87[67:66]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[67:66]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ca6122a (
    .di(al_c665bb87[77:76]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[77:76]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_98537f29 (
    .di(al_c665bb87[75:74]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[75:74]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bde27f0c (
    .di(al_c665bb87[73:72]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[73:72]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e7aa3c82 (
    .di(al_c665bb87[83:82]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[83:82]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_18a068eb (
    .di(al_c665bb87[81:80]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[81:80]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_47c277c9 (
    .di(al_c665bb87[79:78]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[79:78]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_46b6f6cc (
    .di(al_c665bb87[89:88]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[89:88]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7950cad1 (
    .di(al_c665bb87[87:86]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[87:86]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ed72a298 (
    .di(al_c665bb87[85:84]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[85:84]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_49f45a2a (
    .di(al_c665bb87[95:94]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[95:94]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_cefbe42e (
    .di(al_c665bb87[93:92]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[93:92]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_fa2d18c8 (
    .di(al_c665bb87[91:90]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[91:90]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b050f7ba (
    .di(al_c665bb87[101:100]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[101:100]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_64ef40fe (
    .di(al_c665bb87[99:98]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[99:98]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bc89580f (
    .di(al_c665bb87[97:96]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[97:96]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2cc56313 (
    .di(al_c665bb87[107:106]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[107:106]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d3b94c51 (
    .di(al_c665bb87[105:104]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[105:104]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ed66ace (
    .di(al_c665bb87[103:102]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[103:102]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f01d2606 (
    .di(al_c665bb87[113:112]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[113:112]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_61bbe869 (
    .di(al_c665bb87[111:110]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[111:110]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e9846b48 (
    .di(al_c665bb87[109:108]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[109:108]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b919cc83 (
    .di(al_c665bb87[119:118]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[119:118]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_851b239a (
    .di(al_c665bb87[117:116]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[117:116]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d0a3a789 (
    .di(al_c665bb87[115:114]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[115:114]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_db55c0ad (
    .di(al_c665bb87[11:10]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[11:10]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d5c0af67 (
    .di(al_c665bb87[9:8]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[9:8]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_39601473 (
    .di(al_c665bb87[7:6]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[7:6]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_16536f7e (
    .di(al_c665bb87[125:124]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[125:124]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_46fa69cf (
    .di(al_c665bb87[123:122]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[123:122]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9de7d436 (
    .di(al_c665bb87[121:120]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[121:120]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_415c1c42 (
    .di(al_c665bb87[131:130]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[131:130]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f5f2200a (
    .di(al_c665bb87[129:128]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[129:128]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_aa117729 (
    .di(al_c665bb87[127:126]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[127:126]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_44e6e8f9 (
    .di(al_c665bb87[137:136]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[137:136]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3c7742d (
    .di(al_c665bb87[135:134]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[135:134]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_73402ea3 (
    .di(al_c665bb87[133:132]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[133:132]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_26ad8d0d (
    .di(al_c665bb87[143:142]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[143:142]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ff742404 (
    .di(al_c665bb87[141:140]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[141:140]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_792aaf78 (
    .di(al_c665bb87[139:138]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[139:138]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f4c80c53 (
    .di(al_c665bb87[149:148]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[149:148]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_121e13f6 (
    .di(al_c665bb87[147:146]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[147:146]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d3981b67 (
    .di(al_c665bb87[145:144]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[145:144]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c141520 (
    .di(al_c665bb87[155:154]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[155:154]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d83f223f (
    .di(al_c665bb87[153:152]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[153:152]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_66b0d132 (
    .di(al_c665bb87[151:150]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[151:150]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_95ccdf3c (
    .di(al_c665bb87[161:160]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[161:160]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3a6ff90 (
    .di(al_c665bb87[159:158]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[159:158]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_918bf288 (
    .di(al_c665bb87[157:156]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[157:156]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ae15174e (
    .di(al_c665bb87[167:166]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[167:166]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f32244fb (
    .di(al_c665bb87[165:164]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[165:164]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_570f6af3 (
    .di(al_c665bb87[163:162]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[163:162]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9cd9d4e0 (
    .di(al_c665bb87[173:172]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[173:172]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9c8652a9 (
    .di(al_c665bb87[171:170]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[171:170]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f9217ebe (
    .di(al_c665bb87[169:168]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[169:168]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_6a85a0d5 (
    .di(al_c665bb87[179:178]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[179:178]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_fd412834 (
    .di(al_c665bb87[177:176]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[177:176]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c864900c (
    .di(al_c665bb87[175:174]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[175:174]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c17a48e (
    .di(al_c665bb87[17:16]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[17:16]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9d54b17f (
    .di(al_c665bb87[15:14]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[15:14]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_8252cd0b (
    .di(al_c665bb87[13:12]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[13:12]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7363a22f (
    .di(al_c665bb87[185:184]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[185:184]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c73b750b (
    .di(al_c665bb87[183:182]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[183:182]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e6433d11 (
    .di(al_c665bb87[181:180]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[181:180]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d4143cd7 (
    .di(al_c665bb87[191:190]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[191:190]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_cd8197d5 (
    .di(al_c665bb87[189:188]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[189:188]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_227869d1 (
    .di(al_c665bb87[187:186]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[187:186]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b77ed490 (
    .di(al_c665bb87[197:196]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[197:196]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2d5d2050 (
    .di(al_c665bb87[195:194]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[195:194]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ca955108 (
    .di(al_c665bb87[193:192]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[193:192]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bf0a92ad (
    .di(al_c665bb87[203:202]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[203:202]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_a60da97e (
    .di(al_c665bb87[201:200]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[201:200]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c0781ed (
    .di(al_c665bb87[199:198]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[199:198]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_43f7395 (
    .di(al_c665bb87[209:208]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[209:208]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f6128a4 (
    .di(al_c665bb87[207:206]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[207:206]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_72f7da6e (
    .di(al_c665bb87[205:204]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[205:204]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_fb1a0f4e (
    .di(al_c665bb87[215:214]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[215:214]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f8bef5ac (
    .di(al_c665bb87[213:212]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[213:212]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2207ec0b (
    .di(al_c665bb87[211:210]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[211:210]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d16ac154 (
    .di(al_c665bb87[221:220]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[221:220]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_75c0a8cb (
    .di(al_c665bb87[219:218]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[219:218]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ba5736de (
    .di(al_c665bb87[217:216]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[217:216]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c76cb117 (
    .di(al_c665bb87[227:226]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[227:226]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_a1fe2b8 (
    .di(al_c665bb87[225:224]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[225:224]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c7850203 (
    .di(al_c665bb87[223:222]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[223:222]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b4c755e (
    .di(al_c665bb87[233:232]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[233:232]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_669fa2e1 (
    .di(al_c665bb87[231:230]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[231:230]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_a97a7e75 (
    .di(al_c665bb87[229:228]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[229:228]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_5fc18b74 (
    .di(al_c665bb87[239:238]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[239:238]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_37e5bb2f (
    .di(al_c665bb87[237:236]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[237:236]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_f18a3c09 (
    .di(al_c665bb87[235:234]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[235:234]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_240dc3e5 (
    .di(al_c665bb87[23:22]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[23:22]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_40e9c2ac (
    .di(al_c665bb87[21:20]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[21:20]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_809c9756 (
    .di(al_c665bb87[19:18]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[19:18]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_cc42ce76 (
    .di(al_c665bb87[245:244]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[245:244]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_daf67dd5 (
    .di(al_c665bb87[243:242]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[243:242]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_2d08e5a4 (
    .di(al_c665bb87[241:240]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[241:240]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_d0a339be (
    .di(al_c665bb87[251:250]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[251:250]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_83076777 (
    .di(al_c665bb87[249:248]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[249:248]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_dd98c7e1 (
    .di(al_c665bb87[247:246]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[247:246]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3d8fcfe1 (
    .di(al_e8087d79[1:0]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[257:256]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bc848f2e (
    .di(al_c665bb87[255:254]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[255:254]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_bc7c8350 (
    .di(al_c665bb87[253:252]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[253:252]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_954320a7 (
    .di(al_e8087d79[7:6]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[263:262]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c1fb8950 (
    .di(al_e8087d79[5:4]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[261:260]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_62065d1 (
    .di(al_e8087d79[3:2]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[259:258]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3ededa55 (
    .di(al_e8087d79[13:12]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[269:268]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c35be1f8 (
    .di(al_e8087d79[11:10]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[267:266]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_79522b48 (
    .di(al_e8087d79[9:8]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[265:264]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_47621533 (
    .di(al_e8087d79[19:18]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[275:274]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_4e84c1ea (
    .di(al_e8087d79[17:16]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[273:272]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_83909d (
    .di(al_e8087d79[15:14]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[271:270]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9693a471 (
    .di(al_e8087d79[25:24]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[281:280]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_dfedb4f7 (
    .di(al_e8087d79[23:22]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[279:278]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_74e0c78f (
    .di(al_e8087d79[21:20]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[277:276]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_666b9366 (
    .di(al_e8087d79[31:30]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[287:286]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_c9ed8807 (
    .di(al_e8087d79[29:28]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[285:284]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_de814988 (
    .di(al_e8087d79[27:26]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[283:282]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_9ac21e0e (
    .di(al_c665bb87[29:28]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[29:28]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_e46090ab (
    .di(al_c665bb87[27:26]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[27:26]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_cd580b67 (
    .di(al_c665bb87[25:24]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[25:24]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_8155628c (
    .di(al_c665bb87[35:34]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[35:34]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_7a3f7812 (
    .di(al_c665bb87[33:32]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[33:32]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_50f3b778 (
    .di(al_c665bb87[31:30]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[31:30]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_94b2d8e2 (
    .di(al_c665bb87[41:40]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[41:40]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_3e6ae697 (
    .di(al_c665bb87[39:38]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[39:38]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_996f6d88 (
    .di(al_c665bb87[37:36]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[37:36]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_49e7cbd2 (
    .di(al_c665bb87[47:46]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[47:46]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_ec0fb716 (
    .di(al_c665bb87[45:44]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[45:44]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_deb09c45 (
    .di(al_c665bb87[43:42]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[43:42]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_b751122 (
    .di(al_c665bb87[53:52]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[53:52]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_38f2fc04 (
    .di(al_c665bb87[51:50]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[51:50]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_1d9c1b22 (
    .di(al_c665bb87[49:48]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[49:48]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_faa4e9e7 (
    .di(al_c665bb87[59:58]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[59:58]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_6a82697d (
    .di(al_c665bb87[57:56]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[57:56]));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(2),
    .DATA_WIDTH_W(2),
    .FILL_ALL("NONE"),
    .INIT_FILE("dram_w2d32.mif"),
    .READREG("DISABLE"),
    .RESETMODE("SYNC"))
    al_62d3643b (
    .di(al_c665bb87[55:54]),
    .raddr({al_af133298[8:5],1'b0}),
    .rce(1'b0),
    .rclk(1'b0),
    .rrst(1'b0),
    .waddr({al_9c7fabce,al_6c6fd169}),
    .wclk(al_ef3696df[0]),
    .we(al_b03fffe1),
    .rdo(al_8c7bed02[55:54]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_b0f3217d (
    .a(al_c394d21b[0]),
    .o(al_a3f66965[0]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_50ed221a (
    .a(al_c394d21b[1]),
    .b(al_c394d21b[0]),
    .o(al_a3f66965[1]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_6689889a (
    .a(al_c394d21b[1]),
    .b(al_c394d21b[2]),
    .c(al_c394d21b[0]),
    .o(al_a3f66965[2]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    al_8c709c49 (
    .a(al_c394d21b[1]),
    .b(al_c394d21b[2]),
    .c(al_c394d21b[3]),
    .d(al_c394d21b[0]),
    .o(al_a3f66965[3]));

endmodule 

module AL_BUFKEEP
  (
  i,
  o
  );

  input i;
  output o;

  parameter KEEP = "OUT";

  buf al_3b44a3e9 (o, i);

endmodule 

