


module hdmi_edid_wrapper#(
    parameter IIC_SCL_DIV = 125
)(
    input wire       I_clk,
    input wire       I_rst,

    input wire       I_edid_read_trig,
    output wire      O_edid_read_valid,
    output wire[7:0] O_edid_read_data, 
	
    output wire      O_iic_scl,
    inout wire       IO_iic_sda
);


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
paMYjjcG72uBq/MjFhgv+D2KvsP1w6zWySFzuhyX6PhyNnmVK2f9eNd8xQzI2j8J
PpXtqBrtu/Y8QXH0+7Wk8RBQm6RC0prDmA1X7I8qnGXaUee0jJMfvaxiHD6Lldtm
o3KS2vmQq/6P6Ig0+C8lNzWoyNed0x6vH0W5HKkZBpM=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 40256)
`pragma protect data_block
bE11SXp3MVdyOU5UR0N3SrU8mLPS8aJQ9fwAVSB8wkOa7ajOUDvgn+4Jzq5bBMuo
ZYDTbj1Klj8oBFQSLV7RtSBUlWl74+ptE2ijQ+5sDULe3a9/QjlkE705HQTpirJf
lOYVgQSgS2+vPMwyQdrcp4q6l5WrycN4yxFkUT3ilFFsbwadw8yj+duFuYvj0rU8
jdrVy1+UDuPnLE9+XaYGDNjLN6uBoOL1ZljJfHdQ7jRItpq2u8S7Y4fb6ZriKY04
iImPTeFmIfL6CT1LiXfWTwUxUr6AMTfqlhpKW1Ow1gfLs3RrrwGT0tVbw3vX2i8w
X9kGMRLrZJoTjlqOag9b2hEb7DbohWmOt8DN+pmF4qeXSKMfERDLnNcQx6Pbcl0K
06CNgIcpryxo9eM88UPEi4/Hn0cmbQ5Q19diuphLAxvWc64/kDlSXN/dE4VkoiSI
iVVri5fTzuPBXUo1p0eXbD33ehqD6U2vKQzrlw0Nwn1nfSjKJyqQX1mbafzzm7x1
UP07TJ3HUir9ItmIy6o4Ciq7tLgZYzR8i/w1/p7kDr3jcFo9kjVW8RKopoYcJVrZ
bpD/Z06aJJUJWSrLDc9Myf7cmFELxNEaJ/wfYiPjM7SZX2yLuSinynk/BtTG4scH
EozeknPUedS5G4YIRu5AG53paRlp+QO8cbGEJc36MaccdEBAVVo5P6vqk1iAquno
4qqEvorW+YwTckLou0qEsf/j05mT2DJ7tPRox90kUKu1vTmfe0QEjvaWoPOgxB8+
i1fbDBlE9dYGATkhehlZEo6Am3+9eBZiMWxBNlmpCHlRmqcSo7OU+ACxniAtbYAG
GNfWJmrUP/DWXqmQbgFuUzCd3947NAj2S63rAsNArb1FZv5Rr7KO/zzLM/Ah9uO6
m4teMyXJguwVRgXh/1gEybuya/yApqs1X73pwHtp2yJ1V/qVGwU2smueWevoLWRa
2+wyLHVPMuGwne9LhuptvnuVeeEIAKaz96I69bDLJedDG17lXl+DHxduVu1uXay3
n5U/87RW8FNAYdwBCio53Sz6UnjnD7ZGiS7eCMlYC9LYGxB7EVkCOSyiiyfBPuH9
r1slrPEZ+NAZJrAZsZ1qhVTwGnHs/4U/COrlR0rtf9R7uwhBT9bSFsFrMNhFw044
Tjm2frApR8JnTE215Gb7FdFdZ6gOp4boJ3edSyJdkJBfhEVistpvUQYg37NmM13O
pIn1opfNBKhOeNH0433Hjr3Id4GQkKI9G23rVNf7RZAdqU6lTgjezayZ4qIYVGzF
0XyYKn2zekzEdRAGMO6Vqxa64ngQ0c8axytRWWaz2HktbXSuwyikTnQlZ1cSPdqn
+aEU4UyvQlRsQyY4Wqh6K0L3Kiqig3ac7ne1QavTb70MxD8C6fjhoTE46FcLpOfY
EoEvx0Dfl2a5f617Pv/3KQvraD293zqPQ5RZckNWbzj/kld/+Y5h68jIBeBCsTTW
y53i2kS0Mhsc5br4euXW9reJOUKqUkAnHcHZz8UcQtTZGr02xcyu/M8xsPBc2IZH
53VRk5TegAa+TlxS2NlTfC/f2rf2hdmeyilGqVF43/kdEu7PBuNrZIL5kEC3fnRh
OqCk1TL8Ra1bnzU4kWBwTgoZFlZ3yfuf0fTd8MouuDj88NMaTmKa3ErKzPlhJYX6
QSm+SDUJVmlETm+X/QFZ70lMAW4L4Mb7W8LY7DcdrR81Q/SCW3t9EJd991xLp5OO
nPb11fQk+4ndTgYncLhch83eQhOuadCaG+CrNvjMFGY0uJVjFgAFusGO6sjU+//W
mAAMn08FpF7ljGqsbVr+VhyxDKICAleeHknYoXhA/oaz/PtAHMJDYcexpaPA43gy
PveCydeF0C26pP+OcSp5uzHhZR+uvYX54ITwC9eCs/vJWDJpS1qJqSAvyFdna6N/
LA6EJUJqwml+JepgBgN45amZO7ccoaAy0tw21oTH5Ost05ZLl1KCOgi5KZlrFGgp
gSFaiGPeIKUfVWXRUnFZ0mXmM+UMGzcTlkoTDrn4OTvkZAydIHAoboyhONS7chhR
prWWT1++UUh3qoMTX/IOEXOWoQ5mn3kwvAK9Wi+63/ysrxbBPF2cq1cJ82xr5uBP
0zHlnDhzUFB6u4s6rOaQxHAG/oWfOKa+IesiQtErxd1+GRb+pmq2a+GCE8LtSdlu
ERy55BMmoUsXchSBbXAdJ6KmaqMrOfZeU1cSv49bgqDq+HeoEXMkG0/LadK80N+w
S4PCJXwQFpnE0TU+2GeF0WU/LbtvjNZicFWnv14STcHK5H+9QwcVwZrIHmqDGIAZ
KGBHtbaBvFPl5r1jrGCo1WHNky74pGHiRdJtWNUpkSGug0ATYlVRWUnsvw43Iwm+
TQ83kebqSUedwmaU0u6xfspc2P4O/6YqwU0wkJQlQRHjFphzFHsGt8tTohBxWOXJ
/w6nEwLfw/TEeTSAxNIZ0IcR2wMbzVsz0g6uPutUofhmqdiw4q9AW5Hgk7GrJCer
2TBUgQbB/VdDTKgMYf1exAVAfOdrK8DFHQvyYjYho1x9SAvxJqXkTmWG1CIBDh/R
ODQY4gXdrrwxc1N4uatg1f8ZDcYG6rR1crwhs/VWGAGsvtiC43UWsTiEDVoD0SIM
8gMbuC3yOloUEYnWBbTirF9WAkxKTPMQkTHNx/PKBz/GdXkD9bAiUxMtUT2o4svY
B5VGcg9kRH4fl0gGU2Bh3VP5jD2qM/iF/8M0YU63wEdDYVRwgNOZl5/gS+2Dn9pF
l1mIZq0cMxGfNtNnN8ZUeGKTCGD15r9c46ZPCOGVggJm5yF/rlXH74oumt5azlEu
isEgxpQ8RmEL8l5v1orybw/iDtPqG8ChPewQTeftmHCFYx+z35QLP7HcGizB17jF
4/CJlYZSNBVSc2FhK8h1CgiQ+/qFwf+UebHX05bu9S+iKBOlr6SpCULWqyxwKzeF
ge5egY30ySzSudhx6iJ4j+U8xn9FtHQ1a3TNSaRTXANw3Vhwe2EfhsXhy4IdiNwo
BoNw/QmSSJKsVPguVg+K3hsF3fHIboO5joEQJCDFNRWQSGDwZF+CqT2od7WYXLD7
TtV+mCDmCHyOSA837+VXEj3/NGmv3oPgJrj/m6KjVK6slv8WawrBehCROmcdvmFd
k6jCSukO54xvfidOkrqf6Z3wbT7ajpa2Ze6PNBmRPQradeOASWI1cWyqsqexNODD
5kC3LfCir3f51KPhXPL+/FKUIvrR0jEyXAfJtvcEMHed3ZtnZhFHMKg7+bTmhrhK
U0BG/8BFNB3mYG41bGygoCC/LujYCpy6gmtHasWsQTEKRFfWyTO9mO+ZBTiA6o4f
Z5lehzHA4ozYMsitqez+gzArkLT0ivaQfRSs1cBdQYD9y8Yt4NBVSmFJ9vFO9V52
0PvpDHnAs5Ok6DDiVyxmxYsl4gwMElfi1gEUaij2hZ6rG4FU+OPrkBpBzeYi5agI
ZJZblQ59ps8HEnzYv4aPakEC815VEg/+M/xMDH8h7gPe5gqaQsqkCs5UlhkrOyTk
Zby5CF9oHn768BNiT64+pcg16JDTqmDu9INnMZFKx+L6Y49DIT9svhNPaz0NPyzh
G2t0Xng9TZ41YdaoiCuXTZ/U019huFwDz1FoyAlJEo+PbEQM5JS1L22EcgEPGqwL
5/g0CWgNDymYjKXNiFQNcJaofmVhzODcrlKGeCEv23x8A8Dp+ZVv/Lno0DUXuUru
Ip7U0PMdI8aY1r/Zk+SDC7/rV2LKRJ5LL6YKo6T6RvkRv40x8+K0YA58VBETM89n
w7DTHgCMNNshtYqNbGkr3k0mxSIyVKGAU4kK+dCiC7QVrxN9WRqChElph02vwOtw
yv40R3gZzsEJoXB8xOd9gDCZ/5B5uYJEYmNn5crj4Z6axypwqbyXXSQhK9PgDxFj
+FnVQKS+Dm5qzLa2otr9q1RBES1h3YTfeOS51V+SBj+itHiS4uQvUdw3lT6hQ64v
P864mPctMKMZRzH/tzU1+5wcPXxCgbg1fmFgYxKIeTaW5KaFIOvPt99vWL4wZOV6
NAgTbJviG2785TPpZApfKf+UX7WGmeR7G0l4M8rgxbkkfu3Sv7jXIbvMsuI1jrOO
lUN+i6Kf7KBaH0DAXKCGFxfiFMwI4OM2P3n71yEpYMoP/QWJp0viGMQ/1tyDdnvH
v3sB2I9jG1zYT0yRR4cPBeCY4I3Xgt+VYMCCEF3QO+oZ0OoQHHi34qvf0EI0qD91
gCHA5ajLBmBRyC+U6lGSSMfddE7d403JYUdG+cGrvTs81YFc8l9+Flndop7t6mFQ
q6zTZVorJEoiRtkI8rAxX2xz4PQghiPA4dwvQx7162LXDmKqDNO/0etch6PFdbXJ
Ag1INVwcdGUrrFOU9GXjKQDxJkaEW9PahzacVKHV81MZQMXYQj4vOPlUPqwmvbJ2
o7gLmt7IXrhFQarXcHeg/K9kN4/4NvnAWPb0eWca9ZutV2yVP0/gI1sW9Ly8L7So
ZPiD/PPGmbwH4Rljp5BKAa/XUE+GV5K6aZ/+Ykri+CWg7LBFAAAMiZvFbhXY+ErN
pSb0szI0pBFSsKlvOYvasAQMSjYVzsbiEqftdH1HCG/4kXs1PGymiOBLCVvAcLpS
2iO3Xup5M63ugkvarU8ZW11ds1k4/RiADOFPaI+bouygyYDvUxQ2T18WQPgx0W0f
ipuKB8GMNk8Cau8lsrj8rZ1/EE5EiP6WnWaNjp7bVsgEbwggBqIvUYUVJyPBe/LP
/BHVA7xwa+a6WB6qJ2ZDFm+purHnADIHdsK3Z4gjPkHWxYZNzY/HbOsWHVrEaJm1
ismDj+3bovTPEOcGh90ev+fYwA/jzNxaxqEmlOxLLh9G4aU5G+72iMeuvke5UFhE
hEbMaGA3So9eq6nuffGZXVrjCIdNi+iziUMqiTpTM7CKIlgl+PeZ8uN6/YqDxsEb
E+iF9wr4nVHJ2PbjYnYrA8Figwdook+Asl4wsgu6/aNmq9g+esB8Abg8wjF4Ds1o
+vG/yrBfMG3rIKMzNiigM9qO5t7N9gZggCCNwz+OTuBkFFsxidcklVOMd4Fm5QWt
4W+aHhF9TS3whYwj/w+F3z/ohL02k8wnmxyBmUGjYdBNyouvi2pjJS7mzZV78Yx0
/ur5fohykGxF6/2QitTuUSKTboI5BW54x0SU6qutIFc4k/mXWuLEWoSK7/PXOI1N
TxD4q0pPzfgjFVEmq2mANIeR9A+j01R2P/jYuSp9gHOM3jhZ2Khy8RTDvE24a+4O
9zTM5eZBp1w5plNJ1q6g6BnmvqEZuhPqH8ZafQk4ZLKx3pkIa1TomxaahekEF1pQ
eEQ+J81KohCOrUAnLd58Vyxuj6E3cf4mDvuuxwNQnsScBw6N2ARrwYSrO3oIGd1O
A/4pjRwd9X0Mh4KFeVFjPjaKyjupcDIMcRJsI6OAQJIWECahCTJH4D98sO19fgT9
jvjpzbrzvxqzzx0zzP424fkcHtmw/mJ5Tzxf7Br0jxEvK65gKU+RhcQRqMfloBcg
IkcTVHIgYvkv1dPuWYtq63/ojQl2oSyXj3wqH73zb/ANQP7LKzbYPIiVdJa8C4y4
QZMts0C2AUSd1ae2uocFWCa0nu/ZdPghCVSEKbrDD4CYCk9j9LeMYoyL7s27M9Dn
MmFsjXvlfBG2vnagNOs+FvgkZDjmMsHbvNnL4kBK0c/p1zjqvkjkRkUkjaW1na3s
hu3SDK2+kYlbn+luGy1f135mMLjau3MIF7qO3Hbst2VtmOX68p8Gu8brLvpon5Ra
jKmJbXB47wC2WPX6fhX/xuwswvthTYWk+pexspSEcQwOmTaOxj42QgUVPue9Ib35
wC0a7kkzErKJB6GHfvOdbyqn+eGIwyiN8X7vUWP1qDEof9K8KZmdfs44y0K0x2wn
Y84Sg1DPEoXnxO+1VplQcbp6a9rsRvIO2bRWBYKTGofZFMaOMe7UUFHDKBhp9/z+
figBvlbgGikqbBJqknxrpndYBAnACGiD/iInG6TuMiMKI4IO20v6e0KKBdDcZzSA
+n0IZAFUlsJVfOuQD47pimNhzkMYNbzTwFY9KHia7xrfdAn7Psqlj7mDuv/IkN98
VUFsmSZM2zZWQhhPIoeR0s3hLfG5gXmFEBjj6XTqVExSXCUAtk7/rD4ZrrIF8fJ5
iRYmpFntSLH6sGaTy3JAoUttjFGKIll79z7X/gsjUfFMEFA2m4Sj5Ge2dC/KvSeA
0qNsoB972tlES864nyPeeL8jc1O0G2xzZTeEhlni+46e9LHQfiHtOiIwRm2W8uqD
vkzlTxfR7R4qRVZoieV1zx34k94fg5B0SOHw/XzeaaG3ymU3ps1svtPwHspuHV5l
f8SXXz4ymOj+8FLjmJUh5k/kBsjua0m0jvePKBbJ9MDFyTk/l58x29M2DDIODAMu
J+1R7PEtMY5Q3mx2/mQMT5JGSWj3Ycv8lsfP6Jk/YMjINeI2jEZl1T/3vel5EyYX
MMeI7QlWYSMQHSBq5xfHaD96wus5AhQlFPYDaBQUtN9lIbw59ejqZbzOU5stxFG/
l52Tq4IhkHl/+noBD1I1945q5MqBhjFUhyYMAGPHs4YKsE7V9oek5l+BSEl5bZqV
7Kxt40/nEThAi3rp6YTOu6kVtpAiQqPR/yCHqaIgQoSt+9wUwg/yXGkKB5P51wd3
Snaoc4YonCZo4t6slcIRWU3+s32rw+blJhrcm9BQYlSxEF9AZse7wVD96M8x72JU
3Ti7K8tRtK1xDYbZN+h5IXvyO2uABl9lQp8oFSBZXbhVklt1O2tn0/E/QWoftuAo
ItUGULS/2OyZDICziUS0H6I6eMjYhxag+HqIZRkV4lN0wVaDedlgCvJNkhBYnZXd
4SjcW/hNe+lAvKLK6nLjlEAx6rvOB70bC+sK8Xtt7EzWVx7RGUUUHLtqxTsJl5PX
C4SJLV9flofNDNj7W2bMDDtGfUbaxhc3qGCawpWk47mYiWj/k51vpcSfrZwA+/P7
Bq4ZLQBl/CJm6WbMfShi7IdNavJ3kMzkYkQmJbYMnzxwC1AXrrojZtdUEsN0hQSL
pbtaMTasaw9XILlvv12wSrYrnPe7NqwhGDsQ5yJZqBvjJeBlQKz0jo3yBzLoO+3w
RUc06uXDe7DiOu0B+NJmxNGA6QYhxUCW1in+GglWJlI4DsolqXFqf6vFchCF/YrC
5JuRFm1FOFKORMvCtNjpTv9LgnbikBJ3i69ZifWiAWq5VCvi8bQ/HDARiJ9MQmMi
RuD9POqTbp9Az2qMwg12fIgj1s3M7VUx4qHHItvk8qXNUO5y0CbPtfi7/1NHWr14
TR/GJ32hLKdQFWYYF+Zew6DKjaQODowJFFqYN1nEy3S5dkTgu1mtpDgyn5WJ2p5O
HlEFoch1un5aH3+pepY6VBUmYsG0DTxbgcP/7R348dJqwCZOiPTFtUf2L8tMWeUO
iqkbgIbjfR+vPWtWQu2ZLEVG9thwsinO6SCPKVooIfDjs6f0XNINjjAlIni91ZBv
s4RkR2EsLCksQYvvDswQP9BYtZb/r6c34NMlue6PC4CW5+f8On221etCyRXPnZ//
D2dABtJwKX3jrHhsupZdVcz7ZU+7/5F/t26NNhtq8QLdXOllx1Nhm60H9S523T5k
WbWYt2AhRBXs+jRgh7sNNvyfDt2ZGYiS7fIiMdCk3EkcdeY8L+cLRdNOH9mw2VA7
6FaaQ4lM98qA0mmn7UhFNsYdgzqrLdK8Yyj9s0ov5Fi7xnw9H8WxeXmADp5QpJHx
yBWWXXJJ2epuXwKQa6e7sogRM1thratjo/9A8L6QM5mRMiAmz1AXX21LEHDGJVtP
KBe+OzXJO+cGukVVXXKuHTbFen2vCX9wVzSK8IuzPrIT18JchLFEtBGEqBYO0rQx
q3bWkUYoDVeRXGfn86t8u+93FeGjtPABqfyAeTLZ6GOx1+k6hxTDVBSbh4dkOEbO
UBjdxwWQyPnUjdtNcP7Cdu91tNzma67NNFbhBxa7Ho+L3pgYhaH4OxJvU2jJZ1wx
WQVJm1+qs3vtWkAIEmhX8e/ZGbKmTpt9jyDzFj3Ht5mElEBo16sLdlaXGp+Kjju+
yLKeqyII2SIuwArzq5wBAXFCD5uwZ2I39zK2YKOn3jkYUSw9/7aMsooXUea6zDDR
UqIKTDOYLtayti31j7DU1lbVKxMJr/ONWNH269itbtc5hjVXftkM6lelJdFbBq4a
iUz2tYP+OeHtkrKA2CrfdgBYP3+9EGpgY2tkxvR5fU2SmfIXkGz3dFhiBPIvrQIs
czaH7ztGVVRegMEej7xLU7SqNhpJ4T9Hs61Ku3cHZLPmVPcBrSpKjVrF1C/V+ijH
UAaMal+wmNz92wHQ6sCKwr07eM/I/KBFVE9y0riydZkldKZrvm4KMo4wjo/Xfe9M
lXYH+wtn7xJ2KxGqN0YgpDAS2VRp5VypU5NA6wnyFNYmUJvXxTaCmVbeIOee8487
2EIo8HAZFedPDJcYVKFFwoBhULMUoKvKlnoJnMOP/IzvgnRhUB4Ir9O/U+FPO2rI
ZcS80lsXSgrRmoV1Vo+jFjA63ad/6cMOZXtB8mhAnhqXzsVx7RWmo5tzIWkI3UOP
2t/UjLkq7JDJRxJLvyc1q1/YZQkkeMWD7uOchfKQ0KH1zosqkS+TwlYLuRe2cDA0
wc13xGz1MJektBKu5ZempEAU+wRuGId4vSxU8DWfv7n+04JQu2rWqiNFLFFG8SVv
0BrnVepo2oiKiks1WlZAZAgmzJ07pK/Y8rWyTciDDFY5vBC7wgUbxl8aGf+u3KHD
vGadMOeI3+YVzvns1uvmKmyskpBeQAV6jIU5uuHK7MQQfD5CTKxCU37opcPFFMx9
JaNgb2FX00Ccf4iBKXmfT9A+Mze+wn8Kam914u7IEn8NOr1q9Id2deMHAH20hMwm
x3IsX8YVLrfsGCJ1yRaerO1TjM97/TaXJMWDxG43T2DWht7+/lxTv0losWfVnfqa
/Yvzrxf4JDeiQnbtnIw39jeF2YU6M4U2C4Le4srT017ghcEOeN266hS4ph+5Q+4o
ZTBST8iQ79tuTBlHQk728I2C4rDXEibQ1AxbgI9myKkrGmv9Kc6oPIzA9eVxHmTt
fQlxfeHE6X1w5pWSKREm6DBCmUXR+U5UHRlKXUV99rl521+sfFDWopzQRM1BbrFm
F3BB6Rc7/aBQ7otKldWfkDEdRv12nurJFKEX/HzDuxVRggS81A0C49Scn1YSnzGo
tCwenbdsZyOGcEHtZjc7QcGuXalKprAezoKjWXmyJ4bO4114OTMLlryVydHdRjxe
w2tuerVckVkz//7Q1GSeUYWgiERRpWRbmeU9ruUUDqZJl1e/N3VlO2lGvZxLnkj+
LWCiCwCjyTkdV9lqlzSdtOKpcqjssLL/mHxKfqkE3VPl6z+GJcwg6UZ3qsTVcIrW
WmYU/kKCePGw3iYA20ZvDrjx8OoneKEHqe9rDReGTsJgEBFusvguiHWH7Iq/BCnb
aS7UaE54AQGVP13cpEMeke9dwKjPmej+F17f0u1La1jW4+obmV+uaLU8x6IwV3yo
eCd4TGMa+3sPyetoNODyFRcelWwy0xOfhKIPAAP+L2kkwCsjxZkoW2mJPFEEDmKk
1f5UFoXBIdj9vinnZwNDdArEJijtTJvUhQi6pcJW7U+ACCcUEKTQPxJFTgW/NpWo
dFFNosS4e9i3CMRL3YZqcLiVFv+EVScbxCVkSA221xFX6L6KEE7HbsWv9CVAA/Fj
P6sEfl4MPvtKiSPTVdCNoe/O1OFI4ru7YXf3yvq9+HLlq1LXVXdRFQrRppQQvwUn
ZnoXaBk9hmeaP8L3AJ94YwkUEWk0OPnaPyRkI//2C6CMPEwtn/64MLQpdh9BSxg8
VBCll+ZbRonng5CRZ9BK19mKCW3hEQfqQS5uZ5uzmQ95oWQq6RwYGT0rKrN7Hly6
JzOXEcJ7QWI5KrTuK9Sju4+KVUJctqyk6RrKenIiwpOugZfkN+vxuHNjNKAdePFX
+MHeiEGzZOMZECKZeGNV+Gx/JmjwsoIRWOIIixvKUD7oYebl6fUpiDolZjl9/feo
IHtEIWKtuf92to74XFbbkAu++6FJ7c+5VpvhbMmjgBntkjtEdookjD+fmIB9i++t
4Xeb7ANZwOkr4huxwiy5JEJAqPHY/qJ01MbJX+D9jR7DgjV7p1SxPW2AiCMem83G
9cbGtCr/Gri54I75j7olNVkMZIhfUo4W9ky54VOuRQCJctkpO+WC7CUjwFgsVnIU
FlM2nsT/YdbbGRev3PUWBYE56wyGjzCJ9dcRPCO859QXS/JzIK3JaIUr/DcwrtWb
KkJ3bHdeZtOz3U7oS2N7QzGh1HegliS8x/J2+TFioU65htOFw4oLQp869CqMPUtb
50r74MPlOCYLlmIEuTrd9BWV6IG6YAzO4Z63FvFBAdjPsGcHyLJCGIuDPoOFyox3
xn4lfMggODgkYXy1++zAIGmiGzENWhJCnzovoNhduqalOa4ElqmNY8BF/m0EZu7F
7AyG2uh+hwGLkS/rW6A/PwWTHH9Nu8GIOEyp8AqqOU6nE2/aE5RNdfP0SQt0y2bR
KoDkn6bWysjDN998XO/iJ6T8LyLM2eacEHLAoNdB4oYDfB0ptXuqrmin4RbfuDyz
C+iA07L06eKjgDmq8MG50k6JtTfX0VSBXlGpNSgkcw2oV+949IEcuOQAGH8K4B0Y
w2Iuoqa+Z/T1oObGMX7wtT+h1KFDmzMYumw9Cfd4tUxHQp3WU+Yw6uu3dqTo2l0m
8HOICel/bUVIoPBP6V6iBx/YIG4k+nvZmGP24pm62bJ7p4u4hxBZS6wq1SyUUPi6
75WotVRDYQOQlBkouLhcG9io3prPrlQtyq2D1xI95+53fe1dNjdAgvSO84bIDyp8
MKcttxhcgrQMyXXB6GubwsfdZqoOAvLU2a+bT8MReSfjsnzFZzCGH+NgFEMBFU/h
RhOtjVDN8UUdp3kQLYoNJ1XzQDe7gd8tG/Ao6+8f6vgQ6j0H5yGRKcYShSCrXYUM
igC5V+TfcBK8rgMvZnd5NswjXcxxGhTomDxWBIZStdPUqQenJ5p26Z2fq94K8ETG
LgfXB9o37O30mF+Bp0gTHDgxg7/irienEBBKqbMDgbI4yt7zWUiw9yLn1uChPcm0
baVB3Vt6eDJER0MvjDMsWm6ywqQifq7qzWrjYcUOysCmVpM9Qv+6UZy0G43SV0G6
LqkqRivrkBPkZvdwlrdqUmmKMS+MxSnVAO9kMafoEwUqwYCxrgto1UU2brDT8+C/
6pRnOzrK4X0/rgGWfpN1beprYOtv6u7Ejkw/AfIgUnLP5laUUCGzxy28FRxAJxlP
X6TnMuUQVQuzLMm6OaFou0TUk+askmnOwAud6w0Uln5/C1mATTKgYWvYgnj48xqf
Rj9OV2G7QzkhNUjONlqPV/Q3lqSnfpF2Fp++LsuBevLJ0griUbTU/SDPwm/ME1pJ
zZlxtNBbzl0ZH4wfGsJTdGWKO6wYLn2iFOOwA/5A/DurTPalpDei8H5GlnGlaQU6
WF/sITyiUJD2sFd70T2gkJmgTUK0NcVEcNLoF1Qjj7fPGf34ZWlW4IyoUWB2cmIy
5Qx3O13hUfwh45m5iVAtcY8kh35tYlNd/UMHf/G+J4iZDxACVLr4MPwKVET0ZUlg
FyJlbjfzxV6owXJUB4vYYJ/0QExU1oF0aITfWuUwWWxoviaLK8sayywKVq1umAhB
8R8DfCf5ajCGLWQfc2o4dim+4jNf5BX7Y2KH6oobtCZWqlDXhv0O5ds2zYnDR+mu
MFdSgj4pp/Dq2Zyy4K6JgpL0bFX44TWvP8P7Ma13fW4ASa+13UnOW4mAmj7VMpvc
uQCh0f4U6bN8n9cIbwkMjfqG4kDi8LrZpj0WGFH2zW3thGDDa7lFH5xTDYlAw+fC
TcMYw7St6mJ307K9eMpEE32556S6sWypWhATO/hI8iXVAmTY35ejHIKMlzJ/Qmzx
HjnImwKr0j/a4E0wFlzDn2iJs2HbfhaNO/kchWF0hJX+RItT1xzfIkfegDKevi1l
YqZecB6uyItri73n0SRg9ggNkBTmzQidYBs/3/LbR/wScawFh3QyvBlBOkhs7Vz7
2QoShu1Q3YhQFLgZ2lObUQu/6EGGm17NkTsuOwkbyfApWMAjO3DFlQq52VYhuIlY
GzlzPPGXH/KUanHCNxYmcOHenXm9lfM1aQP8b3inPdZE7OJ2Yx+l3CAFLL1w9jEi
mI80NAxvEJEJVeQF0+6XwWpW/6hZtI0eqBb1U5Vo227/CKz4PG3H2gxCsni7JJsG
uMEsj1X1UDgExa/m5Y0Qx7nhje7eFEyRpUyH9llM0TblR9CGS0OjQAZn/AzhTV5K
ruZ2mGwUCE0qIQQtn81l4AcFv+UvHT7kjzgaMduuidROWnvYZdA6eraW1X9yT62K
AMj55DkiY11fcGYqXfczibC0v50KYxOqab2gyEtHiDW8ZqHvYGf49wEL9K6yLVB/
tij4MvIGYPe1ZxjpMV+5NPvkzEnvG+DjlzUFpAAROiYwt9Muxjszs59I6Q0IUFHG
8YG/wiU18fSNPP0AeL3oVSlts8y/aVKBV8LBTIUQMlhUs+7TbM7HrPMhAmrET5rB
+N/bJif/LCCz3YNvAKRRn2lt5VNl7FAmdg1rVNhLonuYaW4UxqW0qmsdmBWJjkgy
kcQpXRO4xrbIF/nstHaoTfbJTw5MGE8O5f7OAJbKdsXKk2UzUeBdotWXfx6B9jx7
aDKOoG49uSORpNvidC8SY9F5mOkUAvNK7zL2FmuESB4tj0x2iDyTmzZkl29EoYl2
pyDW65fsFdOE9Dnq7bGqrS+BD5Myg3XsCoeEs20cQnfH9isLu8FUKJB8ftux1QnH
0BJ1wpicHYconUnVcKy4X0Wki/PY7LEvfiYUQOgwQeW5rUcL6BtC5gymYFIzcza2
e+t4L8ljqvjMSQPIn1zeZJswbG2nv/W/ccITQCK0zqPLYihSJ24Cp2T3k5QZ21wx
zlWFPmk603ljkJKVSGRbWzBBCRCulLgHmNfI//jKtWR8nYEAhM7H4mQZG7ItlUJd
p0fPeR+rXhCHNwS+zUZOBNfjRWUM+kYbXMHDPmkBytzEU0t/cECxXkbtj+H1HF3P
qzZhNSND5qQMDh9PFs4987ftSa9WP5B98AM4ReFDHeL1yF1+mZqogHyZQ29X8ACc
nrphjUb5cx21h6SIP7mLXOSRlhYSQW0QoyV83iOkd4++NZ5ooYPYgA8D81JIQuQy
efb3IXvlT98ObATo7m/cLAGtgVdiA3eoKVrKEEG52gZmISXCgjFIS4PSsN9QOc4d
sYYeAezNqcrhurufcppGef+iGmMdB9XSnzMTA/aHqGwpCMxrWI9ZU6phyCPRs6uY
izu2ngCdty2alRrE1JfItgjzIvw+9/4bzIc/JKM2QUooxoG5SegkPjpYzM8A5/Lc
oqvxKVe5RCcjnIEv6rRRjWOaTK3eRCEVw9pehuQxALDT57nbW6Kt7+coMtCtbyiP
xTx05wjvYqe1RO8OO+n53LQPzSkAbVqdhhcpbC2kXR1eaaK6UMmEox9BuD1m/ZRF
UvFXuTrKxzq0RT4pGfNKeke6ZSMRoArLWxyXEPl6xt5aJkCcHGdKg7NDbLTMYqqM
Zw7tpsJ125OneL63rHE5TnrzPMAvZIrhrYe8CZ7o4IOwaR2YCx0ovVljs/2q6cew
Z9h9kT2xAQbl1CMEG8+qpb6ZrBP/AKehvBZS0YiV2X2wQRRTU9Gw/XEbrbssXqgF
QIFVqMsqgfFRA3Gc01fLFC6qwz5am4+ngSz5nZcc6zF/NP86rFSsS6N6ZAVNb4Mu
sdBOl9vS2RI9G8J10Z4ZPQQ8Ooj0awHE2CJLqvOB9fI21Nzr8ZBsJbtKGy7ZlUvo
hH+iJiPObH76nhu/oAYcuzcOezfnoUWnAn0IWbkxvWzHvEcnMtokW8A0lQtiJs7Z
LYaMoOD1Yq03Zj67eqUw10UoSpxU1dsTEvJkztC/RVViCRZSxv8Wj7FkRQfkTdzy
ZEfyJt19RrtaZIip78qASLNrftgReGFPfFuFZVt2cyprG7vDxrEAztsopJ4zFiw/
JXZwaBXVQHGRWB2WLSpSHCrXO56RItg5hPulSGssHcUKxJ7DQnGd8XGf7Nx4u5qg
ZotQ1VWTgGb7Ic1OT+iaHBbweHWQhh4j3FSwSCIqwm3+qkNMH0WjkigYAQqlU6UI
yt2aFiW3cTk6jZMCZ+m+D7R6l3fbNgKNq04EDaLsCAcCYcK18gfD8Hm3E8Fk2tTM
Y83Jx9ZwByvhfcRzzyf0SDeg/RVG1S2LWZY1R/20kVu8XrRPr6GclKHr7ls9Cyn8
gq5ZJC9NkxgZBif3cni0/CrYCIeAUUWc8WWvfz9XWizCOChenZkrPyfTsS9NGrYk
GI3qIOTQs7XD3++nD6Q5vv5hLa7fP/W7sMWuNa0qxn69NjJDfv75tVF3nVD3M7Sv
g+hMqobxu/35LxEfzOMfo3OCvwS55SrNNhXtmyzHOHWetE8K4BTZ5OSlr+hH+MPW
jrLTi2anRTDXl+P+lnKPrGghQD+PsC6ztlUuxNhx30XWnP26hQsKZWHHnYc5zIRI
B5E+CFw54a5ST1IDU2YL0udqhcxvSTsOPLWwJOTax/sgrS6k+j/SMkoEnm2njGuf
PcJpf1g7JDf2eqKkUN54gHKgpd2+4sr6ZpsZyQA7y+vf3nWjdhTqvO36NjaNLu8x
9Zfi5d7cf6ZOMn6V9Jci7EiludS3kgfZNahRDcW7uJKx/w9NyusYqLBxel5+jZzF
oICDhfZKUGD0EOlPcKwNOaOvlbc9Kf/XCXJ4I6JRVQqkv0Fs4/uPVdxVxf0SFvJO
GfecBwSB69JBXenANMpVYokQt8w7g93eCLcsFdrAdkCdg07/nz1SqJobc98wXatS
sM0xoe25QsGKVfaXDhhVG5yyV3oCSMdlL//M/rv40F7SJ0jPcgLIM4azXTp9I0UH
lBbgv9mZX5G43vQ3suBJKTxhL8EkXI8g7MRBbouHyQaorslvEdB+FGfL4qqpmx9K
zfoOCWkD24/KxMPwu/Wb96uGMumeJ1ZAvGzOkmsbok0kZigBDbV0dStwBAQONdVL
FKjuXpq+oCQk8blIopMvb8tAat6FZMKose5VfVKROLQ/zb2cqlx+kO+UzLImosAS
kwLazKOLgBpLhQCvxsjl5qTc9JeqfGMLns8SlMBsoxY33mWWrOgmbJth0D9fMsHZ
QQeVCVwYkN+YvQmzdb3Y/79IzmqMNlGMvXqOf35Im/bcytkbQSuTrxbGv62hOvqi
zGoGaIHgVdbYwQcaKYU5eQVWMoX/W9fwxDmrX4WrUkSMKylhUSFK10j+/3tsixID
GvSUuYJa2yeLG2GvTkWshdMXSefbFGGq7sB1EyOQ03sujsWqSavjIHzvyeS76HL4
pq3sQPjxvrHkrhPEe/tIsMLGUnVMka4LVBv5T1JjUT4ivzUhljp8WRoO5HBdoj3a
HuPeHDBsE+EC489A+E4oapNV9OWBBOHoMlSyjccGpurXCyYz9kzuNENjNAmWDW/B
BROYUZlEvc24KCxfb9azh1U3ZRAhQR9fNUJ7T6gQzF5saaWFDeLBE1k++aAL4bmI
E9Qx+elM61qLRAYu2CV7yGmZlzix742kphfwjCerI5nQUQJEU+bi/UfOJ9VfU2Sd
O9MddZwwKDK/bDzNvM2wOuVWJuIOyMCXvdWKVmM+ppR926AhWKlDUnw9pI2GGKSU
rBxwiwP6H8F929/rP1w/NUJFhQ2OzbBIeFOcLxfAYlyuqLqSbGzteBp80JvtHanv
jVC8fyM7IKNIWSmvFMX5QrSLyy2tACYulPgsPBE3Y9a9EiA7m4rU/6iw6AcGXS/W
7JfyMCrQHm6AtTaa4J40E3r3LVqpqZ/lpwi7jIPpIX02DX/QyU8zbRqXnzw7jlcS
K1LuKvkF8P78kmSsUFBZHqZLuLWLu+HrYlUucIPw+nCq3IIS18sX8OkXcHPXlqhV
wwZIWCkb0vJ8p/AzmXWFubkYZByee2nbnubke1NuqysMjQjEciNji7DFDRwAAnoY
0XMuAHzn4VHodoQcebUZlwrCqPMNXXWRYr+2BOfgWcoqbJ38EGqWxLISkIoCGa6B
YTKvqiRVyUIpkAQl5opPKE7xx1e8JA1CUKLClrhS2kxasfLJAVnpil3AlTRWU8IK
uBBN4Ipkp9XXK9+I4zOjCgsLKRWC8t1JpkHXq2SQYlfzg0jZvdyYYQnBEmM/Qg4I
98Yka7n0CTBSgcT7K3JKofZOHEV1lOjkaSDuZFCd5oes5QmMNHiZ9gA2ById+En5
HpE5md7ADB8ThD/pwDfa8vw6m9nJNXo70uDQGzrsQqp7r6kY4LcTllyBtPnYhyMm
rzNJO9SukIgvgaSxhxkgwGQvr9vuQo7E5Lp/C1A/YJ81NOrxxRTRiQIT8Sk8CXMf
k3jOoRx8ybFi6kwL1HBsumsqpG4jrOSLRo+tYF6HUQjdJ1XkzH2dOZqPWc7EV/WY
iPtUATKsMSOoSiBUIa6xkCoTIxWbuTWADjjEXzU93Y0MtSrphs/gAz5OoSGcBG4Q
1PWKo4q/wTDpoRRm7berI/xzrllou3KZpYTy+wn4Y0tBjBDqhAjo4lGcBzQBMHH/
EFKYGJRVchlxnDCq3UTOTdp56JlSXBTMGBHCVYhvYOaMz5eNM1YGhHpGR8UtiiQQ
752FlfwC1pCNn+i7+dFgv8LNRqlv0fzfUR6KBcxU/HmYR6o8oqg2MlI7lBi01+hz
J774LmtvanKOwd5nrIYcPAvAC/aIRvnEwKTTmcpW+oGgdF6fMj99UlQwFKCscjRl
YeWwJwU59/GAdqbVeiuqWr1v2QjeC7lw4icyg0b1TtAy7vtsGwTtDZoCa39VFVWZ
+9xboYLa7b6RP1+9Iubr6w8E7DXuD0CiGzdLyZwLfioE1F81COb4ZfuVi8iqHfcb
ymAUyeCR5bPbu43RFkiLuOeBrNz1VbqO7usLcLXwJfiCIDveeNPg8k9trQxIYqOL
81K1iEqW0iGzx8LdwwOTW0pzS9OznECCfoeUr1R8gT6wKgmP2HzatJAqaNOTIt6T
ByCD/bH0dkFP3UKow8mmohNXTBIxg9qN87o8i38KGKjTM4pT2sjYC4ipib00lQlu
M+rFjNOEKHtWG6uxSUzsIoNdFmpKtSPnaLNFnwe2IVENUYEVstlqTao4aSej2ACL
k1hJeKyCQxZ1BeApSZvOOQLnrkSUCmhqg7Ytt8mR1n4eMU4xkeWFimdTJGIeva8t
hAK5cX6tLncTPpr9IdWY3iOB3x0xHnESTHMl1Vg/0JThzRRdPONS+K+S/sauarsD
+R+xNkSJUEN67a/OK4xPg6iyYUF7uJQEfy5B5POPShuJnyDkvAeYkco/UDIhm3A0
87LbbZeRa2T4yd5mHPcJD0Q6Q9n9+IpqBWZaSorXD9lppHPKehXvbRNyY/rtmHDW
BSgR6Qg/3SfY9h++bI/NMB+o43Izcq7ilwMcdEvkIFiS6fJniePJIQfHdI9dc/2N
Ye/LGrcg0YRjVk/XJctNDuSOXscUULRHeewaSOkaPvnLTe7f5b0n/a0XgMHhHJ0W
Pf65avx3DHGnT7WpnxBzh/tjfJM+ipKuhp6JoDVpHYXUItAu3qWITugMc5gZGNgs
o/ov/josAvfn8bm7keD6EIpe6Dyr0GRARe2Yhdgr5GeRORddF3prD+e9h57ejtep
UgFM4172Gy1QAl3zfYpb6IxMX5hwikiwFiS0PbmbvVf5u+1O4XvmTqdMOnLuuCfj
vh7Ux6BSKgjhBc2bE3n1OzkhlSPLm534AojRdkgrKyQ99mZmP5qXzKiybdUTThyu
rZgJ4h2HWzfZoGRenU/Ze4VdaJ5VmELG2cER0Gt6jnlqP3mjnwDTVL+PYABITdAn
D02OskV6gFB73oCvhJt1nH02k9c2I6BL0/KCNw1k88dPW5KojA+eZ6rabMguz7V+
qzl1v4g20mco0ojlQ2BRzFWFcHTNwRNUIu02zW15B/08IJAaDP2F6u1RYKIH/O/g
nk2Qut/MIjNXJHKS8F7udIM6QdbJYeMAPjDpjOxeiYrlpAKT+H5kDBZQXV3SRd+p
SzmPVq80KhGk2z0K1oQWto+U/wUAmEZsnJZ5R0Z3go/MPIqIDFUqeeoDGqEtfpMi
JJLNFUSrGzN2J234KPUfxENX6yfrGb3cNhvjYZ7nTsPrnEiP2gJNk3jX41hMhg8p
Ppa4TU1daIqLzb3El+xIgpLkiMtuzjsq2ZJUqPzTLSiuQaqb0XxGDU21ns4eY38u
Sbio7WcsaUiMDV4FdVqkOsLSVGljJhyw0ct3PVngSPi7et7JLkBEgu5tRKvThUyW
sJjt2XU0La4ChlC4nx6YtuvWL3P5jneWjHy9Hp8zXqfX7gvbFl79IjfmX3+auVPf
bTohqYCdMj/JZ5OSxlSqWI9ZOfU1m2WYteTz2r9mT2HaEElulq6SxxTyEObJdHnQ
k50rrqy+Uhoj6g1hi6tPdviFmVszYhEtnhyXdm/A6YBs/x9WfcpJwM/Aot8gl0Et
r1yOlEL+6Ox8HWTsSFXtYT5yLiMdQZKxJPprO4hSA9m9a3nUiGHKmaUPmbWT7KaM
iMxrdFzRHScW5LdprFhXo00zqlPWnSMDMG+yrRC3uQnhBly21Ex4nVkz63lzOz6v
lKaCXTMnu9vxtiJFUtm6EYc/VUdsHrrUMjW0oW3lJX9cSc0YrJsUMJRNWa4CvF1o
q6jlSMpKIG2miaOoX/W2RixW2AssJ4shaB4YsnlmHP+UkktDUJd0S++FGCFqakeD
obazvl03Z+iLhNWnJvKjtMZaVpadF3y1vqUlBpGnh/1L7FHuCyHm3Ocgd8zIVvWp
xti5RaLX24yWWjj7RXH+fy1Yz+BHmphCcah7BQGW2n1+oD0/cI1HP8R0yJSoD1Fc
XxJwAyWPrPZ3nYK62zSx4xITfcHhWiLmHzYbz10HuzUJYR+33RjVgvMRl3EEVDMF
j5gDV7mKx4uMSSYVxtf2wl30dmxDXIOiL2P0qFKBWnLMqrB9maLKhQGCczJE920h
xwom734Oq+LJMbESsWjl9XZk1ZSOBXlfORN+EPtZ/9hNWgZ0O0/sYOEynY2mMn6I
/VuZO8ydCXs8H+n4CYSL421zAWw5guhUWc234BsCypCpbcY8/2icezKchqBRzWtH
9MhuZYM0P5Z6AoH8Pofr7H14YW08mmkiXyG1RyJzVwSF9apfiru6wgIduqOaxmDD
k75TNRBzGII1N7JMRhx8KRB/vDa18rL/aJLmXGyZBmv7ga8PxJfCEY0nQpSVDsyf
Cj02GuTY17brtNQCPNgyoBrIe3Gfj2DEg+X/VlO6sWMvW9p5OOcjNwpLzXsw0wa6
MbHVdRCC/5VPIynM3Q04vlVZiEZV6DMmqwJyXq4/kAtdI2yvswXd0422XlsdXx8s
wuKxxB7I+HCPOiqE/+JXKBPSehkoF5+i76INHvIo4y3Gb69DYvk1Vp+WiOFTO39f
TWHI+hVl2HjPpfH8v3OyKKkBdDMjp4wS7lR70WevvvIcSiNjEYstYFTaxSEH+Mq/
5UXfCay6pm3bqQsf9GDimB5F7I9Om6O6qYiyfdTflJg4c0OgyrA0gRBdj5F/VTap
z9bSM91MpA02fL21UwVKNxwr+n6NxL3yyYQ0r0H4QcUy2CyBzLcTOICBtVHIAykL
Oy/sW5n79iZymmYSxoAVyPoWAepJn9DNpyjzgwjjIxcpBU5PhZCrBYxkC0uZYtHV
DJOf9UBiPjeSAfHKl7ce+fufmeUEwc6YyCH+ZQZb8wddJzseZaE9Jic01+UM4P+6
Nr8Na1gwJnh2KvcdllpoM+8bJcT9UFJNjITs4tdTY4ICsB0XBJN24h5MZv3APtNk
mUDugKUccwyRMBgPOGQSI2FyWPSPQR2AJJyB7u1bVtjPSakk7dy7p+rwQWlEbB9X
Rt9sg7Mpg9JgsOZwzE/a/Iq+twdd/IoHjtVpOJaQgLozrQJ8eOhvXlQEOr4513uN
J+lxWliWedoUL4G4/8WHijA4MeVkcAsmSFT7IqejJvJumGFx1uiZ682ZhSwH3RME
h+T/qCUqD2VX3eBIWHbH/OmTJLBFVTijRRsoIEOnx1cADHSapKz/Nw1YHWg3koGJ
glGYQYtgmiAe5doBSkrYfljorlNB0GW1BswG8incrk98jyrfLmqXbA+70OXEA0lR
ZcLoQlTRn6vvPyj/qTMHLWwXx6vli5l0Ynxe7Lzzcvb2wFfKO2YSF3dMMs6QUXf+
0+VaAXWSFLjYA1R0Li6Z/IUeaMuwaUCgFZJQG9AsWoq+w8RY5vBNCCbDSOnmSryM
mUuqRIWW4WNMemDEoyyVA+zpP2PflLg9+T91oj3kuQi1v8s/7kVTa5qTBvzuGDYm
HQ9b75lTXgQAxj1wuldQ3g1dVwDljoybgthrjEYcDhk50+6OS+9GYHasyZZpRDNM
oAay4kJZDvJ0FgG3mdOdei6J0cudpYZ6Jv/d4kl4KIhsWWfscxQIRecQeis/SHEm
jdgb+bEpZ4347PWawrgA4q+Q0ECL+ApaCTCSyZskrnFBZOFwM8XkjXNwSfhuKIKi
jcrhcSLV6xZ+oVhFFmW24+44sPMFLEoQIveHilCElfkMB23xRRMsBah+5YLpqyS4
Y4A1w3GVtJwtsPLLQpxWS7y/ZKDZITBBO59isSlyZZCWT758FgD1h3SaUBboMfNR
+p4uqujEghFsakJDZ4Namlf89hIgyTXtyClFXsrFTAEn2oxZ+epCQYiRhnqNEtY3
JWqAZf6/CDJS44PD3NtKZ8IE6tl6XxZ0JpRsjmmQo+IEoUVCK1w+Em2LDuAji/I4
z5yRfEgzR85I8F/Xfn7hvS2nNvHGHcVrBQcA613Of/t+dx4D6WjHugl3NvHsDter
b6SQI9qBF30XSy/VQFTqlh9F7jgkqQYAcdCixB0eCZxPtlIdTUQJt4VztVDkJd5h
oeGem8SauF3ZsA396a1JR3zCqT3sd6BiFjEvi3fzsz/f+u9F8qkelLs2vWhZ1GvM
SObZrZz0lcAa2X8nbF0Rn5KfTJ0LTEzqLur/0VWawkVd/369Gs0lftkAWVHD/54V
3zFhcpeEDmM3XWiGcQArtEBmx+lI8ci93RSuFVGcCP7qVOiveQE+AhAbKiNyFttG
4WcYryT7/PqENxqvu4z7F8TwdAnWdu5fk+o0qCyPMHXvJ80iFX45eYo1lSZKtumY
wEIkFxrbiyMaCexgjZGRW54ZVFVv8QRj1Nn/J0aOy3XJNRUjXonPYW5rbo/XlTm/
dq4FudHu0Ufl1nmrReyuB36HQ8TRLp1g8cUb4xdqexWLpihQy+0ZRCymkh+pzId3
6UL7z55hVbf4kkqQalsV9Ll23C80iSRbS8DpCxUGRUWhgIj8NzfhzNMJPnVetosd
bWF/ewN9Cu96MAbnqTE7z5cA68WdXtlb8RCMXR5E5yZ999wKOdAnhDniQaK0gzAD
4U0+JnFRVyCyooLfz6C9P3JJ2zREUFwjkljJhFUvBnq32GjoQ+d/R5XwY6jlSj2I
+YQWaJRfeUP1Wdx9xw98Yu+NXxXl4glN7mXYLoYOfXE1KU9YntnDO9pPEgOoUgMM
znxdSzFbP9tLxa3M4xuzb8tAMQhew055AOGa2jftL968kNKw0ab6zzPit8zikYQ6
qhsX3WIGKKg+un/y3b5enAT5DMsL8WhjXwd6HvFKmfHkd4k5Bkue1JPY4hgeWWYG
0kteMdxeT1N9KUY8FePdMcjyo29xD50pTSoOmEK5YmspBrrd/4EJdk9S7+runMjU
F8YwkFQlkQxO3vIAWrRaar/39YNl4xrBFR1V73YGv1i4UWr9VddanHtE5G0Yuw9T
Q89v9Yg92UUTzuaIczwar0QCsfmh0FK2nRiRgnP78m63H04H3lM/7ww47R+IpubY
7Moaaokdrrx0PlAU0nO4XYbnMGA/Q1fNPa8LWQXopyxrihlrJqBNPykW+SBqW6fe
9v2tJ3HTP7V1onXc4awNIbg3Lsl1F/y9573M2HnlDb/ylTRz51V2jd6NN5/WKban
Zv0c9G0Qq5T2aQykcgMXNSAEP0kWp7BircCyobkkqUzGFGVRtCtS+lgbNb2WTAIr
Y30ax5/nactyyZpAHOUKkt3jB0UQ5cQUT9tPw2vHqySf924QFAaG0739lzppOgKJ
HFpysY14Un+L4w42IS9+f3Zd2/X+SJTc06bPMC/0FC+LGJ9vVNyHKjH+zKvd0do8
vRSNkzpdSyRzr5z+mHvuFdrKq8w8Hz0hcqD1VrRhMoEQ4UAffxyyFXOzV8hay7ls
IcOeHOmPTO+1gULS5P5qB4CzSPoPP5b/oxPGRmat19b0iXRs+mux79AtOFmZWNTD
AGXJMNtu/EqkZWVET0754D8FcD53TT+qrOjUJ8NXOlOusDgfweZ0ztGrlh9F1YnR
d61kmFTlU9xqlWvGPxsm220C7cvqeW4/+Rc6yjqG8pDE6QQuMwwQjck2Fsi3mCLK
ZnAQ9srOySx7fQyzSDzy+540dx2Da6S3GuDQ5Bv73HiFnnG0n1dXovOfp/PXumw1
eiSn/nWbbmlJ6O36JPPNKZM8JQJ6ZMxI57pBv0AxuzEFNc8+vgt6CoVa2STMiLNt
BhCK6u/EbRrwOemJQg4iUrB3wVIhMXDHWG/IS179Kfs/NvAYIhua8f/XH4znqb/n
Wtel8gbZNx5PlgXoqVQdCDwAh3OVd2hbTGr9HK5Xtkn1IMyx+5jITdrk5UCl2PjV
vIBkkT4C1UeglrsQ2XulRmY2roxDzKBEY7aSdWwrj1zcz3vMtHetcThnoOUUN/9Z
W8oZNXuKyvTfiSUo2hyIiwSwF1vnMFxOVaM1UNFU5nVwsA42R5iShSzi1ZoLteSH
dFtkTv9cMVSNtKRejPHacJNHySSKy1lRRV8cp94zC0Ar4dFbJpKUWjOoGpLZWTzz
RHpsWHetPRcg4DyQkVPhmw3UVcKKjmUSfW94tSi4P3YX5oUzFGLHegt5CoQkCjLP
77JjDczv5o1/VeoeJBxKMS3bxsK31niE1teigFr8jervlkrFXdnOWEvdmFMJ+wHS
JCvH0mv7YiMCL57b4EX5TWtksemRiito5RUbPN9dXg5g43S+w3gKItSK6kjmmAf2
2UMWIoWmnTZhe7mD0t967QH5UtE1aJvn6lQBl62BOI7SWw/WDYPWx+YEPSWQ9EzG
zQQvXi3pDbNJzzUSR5/EMGUwqCCRMWK36dxvk7GoSGym0XudtsQB6JjC/G1McxXP
A2A12mpcZleCeWGOLs8noNICGP5mVprQHbghH1DdtgrY+33AVS0Z7DLOm1WqlUDc
88QFbl1ORhsW8bImf5pSfI1ypP60HrNjYYALwyHZTZCoXr8qAu7DRTHBxmff1K0h
ACU7IUQBpBaCMHVDYS7+FjODIB11QcvnLlTg988fefF6QkgpEIp5pwuj/bizv6Ye
z59Z2pLhfDvRslUhpQl19KhfZQUgwPjR8lK0ZBidN3jabuomf/B9NZgpnYddab9o
ZOYWzj32q8iSay1kZEq5xE5OEnZ0SNSbpOB1l1jwjhKbJ1gBVjcLUa9H6lTXB3z7
v/IQDWatv+HMJDJT0FEk9WMQCZUwv4pEiDs6XWBrsBrXwUb4fOgczUpCJnZkV3DW
/wZuNzrZ7LCEYJkqNPbem/4ae7L477c5baQhTUzi7NqNUey50U8mkT1qSdx8bB6d
o1Jyn1o06cWe3a/Qsek8ESZk4+/EL6BJ8YFEGNdxx95fzuTFjHmn1VAxVgHAhB+u
zVOGzr2/dM2l6mVxRsGB/XTVG+hkPT5NU+RUMIP8nCqR0cEFB2au9t0vzL7nXUSg
4pdKRLSq1TzBbs13Q5fa8g8plJLQxAx4IYeRU6NXSOKamC6vauAB9x7GwrfbLlv3
F6w7Q3hEnrig8iiP3zxI448Od7PHrp9Du/EHmsoMOzlF5ysbSjdYtGlCC9S5T9HE
tiYMO9sV2+4Qy3L0djZ0JVm/uzo7jwWObv9fq7S65pOSgdZqe5n/h8SeGrDj7Z8k
u1XvMio7WQ1FVEdKBjQDb4tx1tjVUGD8SvbKkGNQBLKBSThfd2VzIXKxHwg+CFOJ
a27NLBSgXaJuvdlkq3iPqy82cnrz/VXP3AxNUoHBUnVlb+YZ/ZmEmxtZNy9qX8O3
8CecuaSB8WIWPd1rAEaPlYWF1k6i8qZCph/a9N+454sV0nvu420i2IJIaNyDPWhc
+TYKTRFxP1tcLzK/3hNH1IKFlDwFEPZDCJdL/xxRTt3B598eN+9y+uHRBJ8faXir
KlyXUyc2+2lxK3yvO9ddYXWS32DKV3uB/rH4JBMQWhn0pATXt9n/wRHiKHNPpwoZ
BR6LOFoo7+k75RRv6uyqf0UkbhRmGnJP/3bh6a0gPflEEj2YMHhrU8HCGLl0a3uQ
G7FBzsZl6kf8jXUzEyzYe/PM4t445dDlbsS8bVowNOcBHxDttR+28+JQJmgqUbkO
4H4Glupyx9/XJ4EEcci/Sg/RkGlVsqDKyHljBIG4tYVTHEdz3tldIMR68y69D5cw
ZlvEDA365J624/picp30b+/S5sLJDbIahmSq1fNWIJBiA6QEzc4abcdAjzpBHrrE
3zLEajrhj2C5q5OcsIqFSeAo+3RN67DWa/08hH7zwI5yMpimyUaTkXU3aQpie8BK
IPifLG0fE8lc5Z3VwhFQQKVGpJkh2SlfKrfJm81qsNN3jjIWLVhhnw7+nAQNb9s8
d23y3SpZvngbciIU1luCKCL2cG/wWrHvWn5w/0F7PfIg1NSQfxMhT+Jtns7utp4g
sN/bhQXUXiZ7rZ9TqVb9YZR0oiGvwiLIilwT41RFBhRyjqzPoKd0+rXvgO6FaP+3
fPqo7t8IwA9VDsF6C+z2SYgA6PQpcE+lDnzngrRZds4SYaqLg3HkrZ6owfHxOtc1
7gZMCjRpOGVySfeTS7msdyaONzys22f0OW4fcyXrZaPp+OxKvVG9GSIPRF6ApeEe
HmsEBZm9vkDPmr2TrpL5bE5nm6l6pqeMJsagTGjli5onT8NPJMeQIp+pk2ipPFMc
Iy6yl8Zf33Yebzx15NeKUxoytj7dbzJtivzzdJFaf8CtQzO+GRdnLqPBe5BYZsxN
D4Plb1AS1AqEINCUSSP8siGQh2xQKqpxARd6ya0U8owly0Sftfc/OUONi6ecFSXy
GscrK4CXJiRQVe9Z+alPzPUW/JJsRlSCBw57xQQKBrQvO8eGKWa+4K//QBqmaGFC
a9SECYWHpHCcYM9313SliL6hLYCwDzJNLwhBMrZnMg6PSgbb8UmDicEhynNRZle9
QCTZ5lFWw1hux5Hup2bETL9Ocy2SKywFHc+Vb2kA+QTD1fy2XU/m4sGLUJqIg2Rm
yauD+nMo1Kd2gGgc/gEIwWMsknDKyBhLfbolvNJD8+7YKu5WFDSH+DNLx2NTf4Dj
613QPVEN730CeOfYL41NDCBmCiPp6+2hO8CXeu/g8BS0Zzw7hwwHXWmpC4Ty2Agy
H/QbIIch6BIr7BYRDrNRsRV/m9aZ83xc1C6BTOwfuJxLuRRexaTBhHht0fkdg5z1
FkiNBDE04fLAhkCdepsb6lj5RUTZV3cRqH/iXiz3I0XV1W9+UVJYrf2E0SgSqmKG
1vCFBYBnzgK/blEUhkLsoV1Ke+7DXterFy95YWHsrR58BJenmTMAyciRzD//A7/v
gx8h+33JTwbXosJnhVMWpOmXZlnk7XMV6F9egURBhmmoPxVQlW5pfDwGqt8YCmLA
w1BbadaO1XE+fgJsM/Z1eahE+OtFerpgtXUmAfvpr7yqJ8FcRnaVoSWLzWKe5A71
E+ikxQ8uweW23+wACjyJBBC8wxCHyIuZj/ZSy1MtkDbpzubtajHPQ4tRlvZwPp7t
I/ZJonmq2NTJJ5wmtiVWkhrkKjghaDVXso3qAlRYyrk9HPvktbJjxXnx4DoU1LjL
YIkqnXgt/YzHagZR/zN6hw+qYbnjWmsZy+hEP/cLu71khIf4tAC40TzQNHOmRwhb
3i1Kx5owDRsgHk47kE3Rucm+X7foLyuFN7St6LVvInQY45LzvWapUWrZz/mBfimk
rzsaakzL0L2xWr4x6j9MeAP7LdlnImPUvpRPUelftGhEyvo5pRnUij2khZQnMl2q
JQINQd3PS6rwKHhxhRoLcwOIZZ0JzVP6hAD1h/i5jF8ni7lTEZFvd3V8XnBdK5C0
4UrOtyrBaCAqslda4LPUrctS0IZv6wevPDyEztezuV1M5LtuHvMWctinsscfrcvi
37KQdUqIsCu+HbCupRlm5nJSggVNZS+JOSsb0Xmoj6r4SpcqcW95swh/zHMuzYmV
4AurJeMt3716pwtkZG2EcoAmmiPckFBc5KA24AhmL8h2mbuIn3I2ugqp2JlfRfIW
unkFJZ0Ib7oIMZWR1hQ74c7jzb2IY5IetMnP/06agLw9x8n8CuWXvfZl2AL5bK+y
spqtQVhhy3qG8qACL5X68RV6+lk+qT0zj8GmdwMn2jQOl9TYoNPDhU/fluNFtMAf
cDZCjiRpi/8Q7Rn3hy7pmfdYKbDM41jxrzaEjv/JNrDhnoA6nuQbdKU/ASGCkwU/
Czx+5ywESRr44ipPB4Aprjec1D8N70iGzDNwbnrjyajH7/Qjg/kaBoCBcow+82Ua
vI0eIkEIsLcVlyFJh6nC4g58W/HKT36YSbkkb9r7DHKcQKbQOUyg7EMFE9g1mEfL
OWtG+P02zPi8/M3brE/RCZ2l6zysDLlrWEB5Nzra1nnPrT9uzvUXppL5w6HcelAX
Nkl7IBrRjxUTSlNZjuxx8nIwM46oNNOf4+vPvNjMd5GyUBttzk4MpSoKv/YhvBfS
GV6K2jgLdOLXbKuFh6XnU91tlFyAI0yinYVIGfnKaox/m03DnoNfNr/XZlMX4Gs4
wltu6S/4s8KjrXJqbY2ak5NHshPvDC+Y3VX67nCrtP5peULb3jb1owVdJsbfqL0c
9sPcaAGen3lQIzxs6smpBrkzFMIC1Mveu3xx8yqcpkectMFPhcUpknePdkxj5KhK
8DUoju57q3kkotpU3KfPflL2/srjmjSjltH5XjXUmK2ydu5f3AKPrNma76X8zbqi
TxG/9kPu/e0VjVvHK+VHFNf8dqHp5wZmnqImY6RnOXcDxxdpIA+S73XL93396Ec6
ShZrDvsH/ZBoAqukdJXX4qrH81ASoBqLos3/1eF9eH+U30oB4XKPF8qJuezd1n3i
EBAIG4bCTMkK+HUwvMXd47Lgeh8/WAQt9lkVXv86qD8pI9YeBifwvqejaU4ST7P6
F3kvCEkL2AZIyv8QQ0QEI5e7Is15virhqEuNYPYnsv3SMQA7s16N4qJm50eZv0zw
l8hM/tw5yKsyXA0HZbjytHk358h/Fcx/zTzn2Qx6tQ+1RV1ysXYU9g7LXNqaSAlO
HuqghwQntPpATDePq92MC/9+G0vxkaXAH+gu1qGn2KcHlteVpdXtleunypbRhJj7
uhYSt8GUkE3TfmndhGRTCTdsq1RUg28CKRXj1unKZwJ1TdTQBIU9eRm0jCXDxmIs
xNmayCrTEZioa7inV8CAyaB2s5155LssEhrsjjGSetJ+VEISKUDqMleL+SsgPAQE
wtFrFELSsyuVVlyTUxAFBTL3CLmNDscPl0N/pBsAvfSkPyENVhMAaK1DZ3BDTN0o
4XZ8K8DClACZr5E1DSTKXjP2xlqVI/hxvIkpAUcDEe79PBnCuaQ/K/DXH8sDdMKU
PH7R7uQ97Pc3cetnKuGKJB1DcNvRhKELu3mnSqjHFICSY/Xz67KBdFyR/SJ6dtNS
ztd2631KeCbOJC5U1tFaqUKicq6zHG4dCxejo7zwyUJTC2KAIDeUQ174eVp8frZl
DluBDrwFJYNir5vcs5LiRHgnWNHfdqhiph0AvVCfyjcFDMC4hHB0BJnM3eRBegMn
TiudZNKT4slI7VvDEBhBqOkgxcyU8/bRNBPiEoncvunnyrsXH+c4sqOmzzDnXnBp
HYYX++epayhgl6D1IMtS0z1YKGIYR/nVSyDHaC8IEN6isholRWpIy1VZo5wipY0A
SF0t4jXNRbL1+g9HvsHYkZzGC8N/TPly35xwZsc2xP6+HFTM5jIeh+Pfqnhk8I66
hZa9kTQ/xdDcI5QT22wdAjxFb4lLHauG/dqEsIa/eOT/Z8Dw6VwgzDWyfRcVsCef
RQqGP2Ju/h8iNNdhMHC24OYDanCp3HkmbkNtdnDUvREemz7EJ69Jkw5apBSgEt8G
4AVpQFj7+KaUs/8+3aPtimj7fadZe5lzIE6LNv2W6AT3PSFR8fp2g+fiU6yntGOf
YyQ4Ver5f32tynTlXpTnuLALSjfS1uvv8K8eQLiUGyJf71LIWdglwI/CTm5iy3dl
62wxLS+y0hC4XpFBEGiqtHbZ9qQIS3o7bA0vKxLjYiqf2WgildGqCq7BRt3kTPvh
lYmVtI4Oe7jcWSfpnJSrBgGJV4+DilM2SUolC1WOTSmCLZpXynJw/W/L/T4RKZ17
DM4HJG3rUg4yLpFnaxDiTBKe/F1Ow2XdiU2s+PSbhf5eHbyxdNzP79dqs8WYOdZW
YjO5C7siPhhIp0C3rnsM5h7Wze3r0ErwEp0SFQ1cuROMMq0kMgvRBvvbKrpn6kjp
ii8crBlivYiivDg3/Repj+dOrYnLLs8M5t+hSo/45gA9Kmf/ECl6EkoZATXb28eV
fr5oHpFkeRMoEO1/SuW/A5/nwW2D5l4Qkb3TF7JoHs1PiCr+geja693Rlf/24ZER
2k+2cjvga+499N4FF+h44U3qorFzqLoTZO40jCENk8rUbH0G9fW0ghQM2hwPI9CJ
tVe4Avs62jxGJQzr+HhTh8Br7czSUUt2saGnbh8bulA4IC2DCNXhgNWoO+EmNlht
oYjzkJ42yYOzbhAxPwQj1otilmITwa5EImWqTHSN2bvxTkxJ5O3TF0so5976UrSZ
B3x+L73oESJYh27D3TljqBq9uj7dhlfno4IAco+2G6pSdQsDUfUQZqlO+ayfi04p
SJiGMDMS9/NG2HvNoatJW6imb1jtC5YZQVl7s40NUi3VHzLPS6Tkf0tN0UmtjsLQ
iZ8kiPrEoXcqTWpoW3CkTyCaqsVsl9MOdAKRv51+zPIY914b5yPdgjNMhidDCQqg
vgTaDyUakPczurDGie2qRMZs0NG6q1zIR50DS7uqxi+gRFEumPqE+5NhipSy6MOu
RsfQI44JL3KDP7GYijSj9TQfnIgY5j+xRnSxf5Xk/3RC3oI8vzspfHWVneIuqPvz
c8g3+CQ4oy/DkB24R6me91mdyVnd0CwVfTpog44xmoGj705jug3hx16dLf7rjvo4
C9BsgtTtlXHWj77P5+yDgHKlQFd1XBFWJaYe4ovO3xdwC5QxjkY4iYgrSINtHr9V
6fPc4Es45jaOmgPDVey7zydTV++z+sFSewv5KYuQUCKoC+4wjYwEAx1yazkxJgWh
58qQX8QMOj+C3JV+bxBdxRWY0/4YR67wlgSAV/inyoc4r+J+zHhRs0+0FIAPsS0m
WRoVABw9JG/zwbThvzVB5HK03u6QwjnhzaS3Sviz3VQ+0ypZwEtDQRayp1AeE28R
SwukKJIMBzTScc/zNPU84KrAB1iyXFAkVQZMYQvgjJYOgaHi769zGuz47pK3WmS6
iHJBiWN/5ncZA43OUYhp324E26X+51X3jAa5eZxe3xOjtZkBi0GACXqWmxhX1u/o
nP8LWX8Jl6160ELnfAEfxZqEcGEAPRgwO+jViHZRa+oJSwmrK1AimroXYKyMr1OA
gbRHarZYtlqcMh9toSXqFkOxGaxm50FROIrWTGG3vLvMdds2YVgm94UrL1zPHW/C
J+anE5Jn2fmYipNaSHuDdeKKScP+0QAJajNBxqRtjuja2iLR8JlgPWAhmYuksdK2
Wxbw4j13bEDtE6sQNX5xDhnUyxnTTDm4Y2gK1wni8Qt49sogr9OpMmW7NZrNfO3O
nwwvG8HzsxCox8l2wU7Epk4xzgzdV/tiL0BWMz3gnNLyCHkS5/CFGfjEioPDQ/f7
zTxeFR0T6cRwVa/SZPlfvx+EQv63NT9h5Y6GExEe8NYdxkSca5mwYFMHhEnQ5dIk
rYnZ0Rf61qVMMRIo0Sp1453X07JlXMiMNDwdYFw2dLe1O+VozEWnOo0l2kDZJoBU
uDaMom4PakKZs67/Q9upNcNDtAO3pCWv3OT+DnaODDENi7PDfLi3LfMxc5uIhqvl
LRolLJ7I+FBawQSP3A9tI9Zd+fKZNG+3vPXU6F3RHJj8zhCBF2wD296kE1Odkf8F
eBr3H2yFTgGxq/r9OXdnFB1IQGCK4M3r0NEwWlWxGAMUDxliBckEmSbd5MNqhFA5
Zg3UP5U2Zm7xb0GIHm5ZA3txoVezLi98LMCtxwFERtciP9+XmcmvWl4gyUJinEJJ
MuhxBEUup6Ns0x4LosDfCHvUnhMhBMnX5K5i3a9RgSguMeXcBB8pPOh//yuVxcPx
cMyNaRq5NRp+dQRjyqvO1hTeEDJt3Z2/wNQCGBx3U20uDBtadeErDwFxRL0jd+YF
Itc51O+qsjTaTiTIhZHfdBVgcr21zZkpfk+GlHsEMpPRBD938GAM1h/vBLTF1oZN
xjx/i6L4/F22qgINqBW4DiriF3o2uY5nQDfWlFCNRMIKSw+TkoMOGjb3FpjqnNSu
cEWYwB4JoJQ7j/wxP6qI0OwGTAeKod+Ug5gWCpprHe6HNGoiYXymlYM8r18DmjCr
sSdcG0eAHv8PN1ZnvySVWD/VzHdq8wtVyUqBcQC5wXOiivE1XU6yU2rC3g6BXFrS
P8uGymwPloCsQxkyG1ArHDYJqJ+2fDeTDELQI9CRPwiuUIRIT7R1G/8C8IyeNaGY
llQH6dDyHvdvb/t95Vx3B06Sgx7FEJDU+kYJYqqJOpvAoK7l+YQ0AYSrQzV6n7Xa
0OZPaQzkHmqPR17MeYT2ccZyyUShuLuoTR+ATq5DRaikI/HrMZ3QniJleDC/exdI
5MIViH3Lq/SPlg7gl3PgV0GLGM2HospsaIzwWyeVG4PEy2THHkykL9Kkv9dscrvq
6QqvX7muvmFVKFuRJCn12rm5Ca9NEUXK0sTkoyvJhs82gu2OhtP0NvcBnFDU09Sn
CkRhIR0mVhAZ/uxQuqT2ChkViCetVpoMdP3GpKVIBmuWC5+3FEmYGXRNRKwBu7Pn
lp+PUqnSyUift6IYuPyaMYvCbsXnktjaBoLg9uxYCaA6b+tNWk77IYVJBt/dNUED
wtaroxjBT2S9y+WmiRcyd8xwagcHkyf39jE2ukouAK8rfwyUAeBxqP8XXwMwno06
E1bk1ISIXH1BUNoVFJyL3wdWz7qPXXPPkEPRbKcCrTfk7dds1+kUzor+XLJ6v/A9
YqYV6A+xdy80HiT3w3srN2ZSyNmWzxp9UZJY8CUXsdt5J3Hz+9EIjgcx6v275atc
SrQT584arBo7EbPkIqeWyKKMxuUI62kWvz2tSOjEiiXWvwCJlDEGG6fOhjFdMvYZ
PC1J+Bx4rBpN+X9V4+1waK/+EOFEPIFvk9yb+Q4JqtjgcGn+fQs1xgwlv/dchqdO
FKGXYVe8qz+thi54flWBN/Jm6Byjj88jHP3NQKwkuGMU3ZXpecYjPszRb5Q/5ZLD
6c7fPbT5IHAMgAWLzhAJ97tRKlwf6piy/5alybm15WdtKJAUixGY21SfuY+OfFSr
20YOd8bpxHbnF1e+0UYap3/x3a4gJ2KapV3qZTQr8FHfBNNORYL0y/1mbufWfHCR
ttKxONrMox1njoyGeWZ2aTy1zrR9T9dK6XAZejTeD8WcmCmoQwFCHq/zfBCGGLzc
6NZMTwayxUAaDLVkwJQoij2YfnnzM58Pn01OcFwpYGY/ziJ2G4CcOuOtjux82TsY
wM/bNLSVQlOn+GFW7wPbrtL+IPQtht3rd+QpGo993EhVXc0y+x3e+JhlKLIYA0aT
wtRzB2uM9CFFUhwtZyBXaprXbHRpEoalFghOLiKmnG2MTOj9HkGSqap9hc+pIyAk
XYQQ25YVXQNJRqUuGN0ZXGQwwUT8FRdNbgi3Kup9nH4zxBjGzkWkz8k0ZJmEHIEB
Aioe4uMUvMlnqdfOAyjfDo8rV8Neb+ZfQcf5lL2Wk0ACnSOcnavWdyPmZ40tO/id
Dta3luGQLz2EsVg8WZ0oV2Nb6PKcMAKvH09FTWW0D4XdSKcUCO0tH5pujwSGWs/L
rHXJrA918oc65qUPsdzqSK55PplTBGor+BJJkhlzqHI65qD97Hl3Fm93tN5YxKfU
rVioIBCOoxGO/74ohDjSR71gwZb/O6UOMGaVMUPgfkuQUZdz9s5nFnkusU+XQ3VC
sxzy/8pjQdNP429QVTl85NQPh9IWZcXeVKWINND8PlzMc0xEOfHHY4RQ1Q6ufwu8
pV+W2w1NsbldBofKzinRGLNDyuxEgInPfp58EcZtvWaTm3T6if2dYVU3W13q3FnF
MUrx1Y7fS8V554chK/5m7WoF961NJjW0PTs7QE/W3tvM5VVC2I7OcqSeYASqp3IN
9+4ddZMX/mbfGAZ9PGmtnnyYCA/kuwG0iYqtH2uXwU/I+NJ41CrMxHXQFotHrvk+
FCoMBv4BKA8s2Gv6xu0cu7d0C0EtN2YV56LQjdxltCZNfZBPJYFtlKTMkVcgO5p9
2ZEQQ5hPLEsUlSbUVhoccla1Jo7KvsP2OTaxY5XCq1l/zCD9fKfNUggvQZYkedC6
Y2YClRHqVVI+YKz0aTj7hB+MjWhywYv0z+ysEK7rtgRl6fznK0zfMKRSNkzJUDip
4s54w4beCQ4nuYQkTLueInYHWnfP6lUeKcy6nVyQtUREqcXzVn75FE4iNWvPTNuP
1SgDj6Z3UzgmdjZqIpA9gMUJIO6b+hsE54njcMOYAMJvyzUgUUVhrRSbiq0Pivrc
sD0hpjoG6NFVZ4aIYttDp8EWswVJkMUZSYT2SfPn/UtmYXQ/Bnds8J6mcDajrbfY
AwB6HM86h9bodye/SnSFtLxbtikYA5XS/+vozj+F7EOmUfXGTGbO9fhg5kx5Lo4y
WFO1Eo4ufqT0yCfIFixfF3QjKD8WkrOlP3De1bosNde9Vq1KWrTLU42vLnugTDLO
2MICgLGM+72VcpL6UypU4Jv7QpuxJacW9VgRupF9MjKf63y8N/fipUd3u9Yh6xHN
urbr/OE/Xb/eOwuKxqfsWAjm7aymd3MTL2k8WWAjjgPGeF6dyMVoRkXu6VwCoyX9
l+gpNRI82fE9FbZh90vqAa6ONS3FpTYGRqbpuLEGMPp8aRCXlZqkajnK355jHvJG
+lDYX2ipYa8eapW75ga6sU7cFdxD2XmKADvsx9tJ6nVytZqTPBjUCKKXTlP1HIU4
H4KjdFBXxjzAyoHLRVnzZDJ1i0QVHnxqRXirqLbe6Be8N9hekiLWslk1apEAD4G+
wMLDzeKKJObcshjXz/x7PA4rbX+9ipC7H1zGsV/h2cF/maF3bT3uSq3bbHaBVeg1
o/udoNItC8+h6R3MU6Fd5C+y0tqMh8KNTq3KcWc09Ne+MnNlFicp58jOoPM7fH2a
q5Ykxh0o0Ch584Wl/PMA2pDUWyHyQR1mYKWRKrsyYyW1cvOdML7/El0r6RVPP+Ye
HfMl/iGfTTnQzKeOVRH72AJyRnc9GA+VGzjzPSdxgSx7MRwi6Y8zJ4vgCXEwjpnD
Oc/UVTFTusJLsCscuz3MrCjaFkP8AgrbFsalTbvgJITuN/anKAqXcG7Xq3Q44SEV
g+EY5hYkQR0T/Kst1wZqXwSmefHK6/SGJfABA54srpbvekLWi4aPMKDjAgYslleX
I1AKCsdFtKaMZ+kYY4fJz/zvd011YqGSv/deNqpixlKqgVexXCqBTlEyghQvH4Jp
Rs5tD65fEAkLGeW3XR+2yrWBSlZwO5SbwbhyzncMpLfrFB35n6g7b/TcOaqyP30T
qBGY7NKksYkq42lyxAw2uhiNOvMmkOKp+f7e8ZUJUvF3em4khLqHaPZKU2FoEPQF
YHUOa01fcsrVt1KRXAo1FtZgp1nYSXC5KEb3AJ0dsYzgXdQDjmex85uccHfGmDtb
gAt4G6TZeOWYJhWbfJ96n3X78Co135p+tFXYhEUjJePI/LteJFSGb5TY6JA+pYSH
oBfOrtZjiOsfI3yC77mEFhlLs69SRkrsb6RTZvNrlsCTDPaWJXAkbhP9pr/X4ceI
uuGz7jcqVujouJPSsRN+ZLRIhqKfbcHrtVR5kNIKttcw4sCS0oius6LSKcY2Mcou
RW+mwBaaSFl3TmqK80bPXpBsQqjUBB+xeUNSXtayOLrOTi1PIjBBDM+j1ePeRVc8
P1xLBJuPlh6KGfaaDRKqoW2uPBDsY66XUddB0nZBTOAMhiK+2B72yn0btdLKIHjH
Vcj9/GD8aJq2ZZ0i//umKJXOWOzeOEeV6oxPi0WI906+SXfoNmLMxerbve/zpys7
s44hfq9nu/EtB4wy/tfNBE/RiX4P6rVHvCv4AElYO3d17Vy5mP6wlJWY/GL4G5+H
muUqWBs5sGoc4SWq/NIQXxvdKzU65EMooAGkpIRRyf+iKI1rBUpeWBbndsJVG4px
Xb4qQMimS19ZoaL8WRw5h/d/e53tBt9wMg2ApnqufFz0QiLQdk6SW2zWLNDWVmCK
gS45bWvyfblkBxX0Gd1pfwhZzEt/7DikpwYdaoBX9f5JE/297akiSrkXdF1cnsis
kFtJjfmt60twIcPDfhA/VSiPIvjvAR8OUNW+13DbUAc2rOgbbg9olHgAL/ymJehA
8ocj1jrwJts3vIgh5UAMibyUrht0aZCvN34iTBpQWuTaqRFx8okQipnInLUOv0VQ
RbNLm3AhWZ3Ry+xrSIe5MoodWX6Uh8CfCubyHIdEraEfNaxqO4mC6do2Dc2DsiXh
8WzFioMeaNLbArZuLlXl8nTqTd9V4WJ8MYknt/0a+8UW3ySMNig1Iz+9tu4sTIUM
dSXDmqR2o5tKZLgmmOLnpbNoSV0P9DOuTWPpE4GTDTdlhwwK1tnqIlGet8Y30G4I
qy4Lp4NSasLcAcRBuZXS+D++jww7TXCUwzf2jfWcw6bMvYErk684wIrGgFRzIGHD
ZOIzWwdY0e4KxSvaxd/2DeggUjopHZu2gYcLdQSzeWnUJBlwlEWq3km+88xBe7z3
7ozZgPlaPzvdrBLwCsdxP0nF0tQGO+kjr6x3QHIgu3O/thUIDkKw7RcQM1KmKyxZ
O11aVl4W7xdJevazEg3x81MCV1p9weauHXZ9HYdkorGLZ5FVnpTvYsrPHHSvY76m
MPedn+N/3NDYm69K6PjyeCEOmyNNfbNQYvTo7Wr8ojVICdG5eiPDijpRPxwljsqk
AyOd3P4pzjRpyuXURlRBsO9Gbibfe9yLc+0lzfES1HlmGfUCe7XEkXMLLUuoWV9d
a6LwZ8WaqZSgL5/SpiLBOCKHQyql08SjzRb1rbIDOVjn8px32QfE8XwD4FF/YSvu
F+afBNJhQ+8WYhdCsg9vmPsYDegVvY7yNNr1gQd7xXVuvgZDoxmcUIxGPt90RSEY
O6QnuA6/xW28eIQMWVyDO3qpSifzXfFkMSQmbr8/F3T6eg/iZjWSHVNb3RlXoN1I
Y2NdYDP0JjxfreLv+UbDIXT1NkUHx7E616rHkii/xlry0qISYoYqjwO7vPBiGQDU
CP7OuTIe2k7fadVnPxFlIYMCVZ2UJ8oMGABgwzp/RiNL6zzO84RjJlmfU101qiER
tDYwLibuKgMREFtq32suvp7MUe/bWOaByfmfpfwm/xDSjlYBq8oBaKM0lBz/Mk6I
G9zQ9J0ZpzX8RaZ+AufjI+9yzmeZbwXU376TkiStitvuI4RXLgS4QHoxPStdb5ja
sgBdVjjAbfeNjRvB4UjglneWoJnLZ5hl4UBHH6YYBB7xqCtcT+PfCqgGgXbdIsxV
79E9VdPkJKVYvyE3qrBUze2fTm7deyXfQIJfsVyCmH8UwoogFmH2gfKPot/YHJOS
5mlgDLqr1lk//Xw+TuJ1Yp8jSWxHc59Wq042N2vefY9qfdmUKnuFvLhB4Vjv1qMS
MVJyuREBVIxBkCwUVYeFqlMKOZHlWmJ+/HLfDc2Ojla/2lOEpV+wGqOt9CwewCKI
RNLKAVpm0ercAeU2du0h20J10jcm0xPq2e86AASD1vTrLcuRj69GnF8CFRXUpnbk
AO7a4no/vUSBnAdAWInHEJ8vKWMkoOzc3rLj3Y652PjnDP2KI2POqsyvHfB3zFoA
Eo4hg4KXffs1FSp1QyNvJbWMCXpv00Aw51OiyiF1JPjtmuzOELq40fmgzmYBXmSX
nqXwv6RjDeCxgwZzwo/iSywsiyrtfQ8rc5/vkGkM2b0ojAQtZrVcPCJilsrKnlCi
RS8DYDGmX2GCxmzBEL72Z/3jzTI6/3lfN8vKY+IUfhrAA9yWHfjzng2f4YdL5e/U
8A1AIt/9Q1B9HJmkPFNky/2mXi/irIcDPD7rzYSoZtcki+M+NeZh7ScYKrErzQ2c
vtQo70yZfnPrg3txw85Mkj+AhrlCVJt45ufcl6pFjl3lg9cDwxpqv2n/fH+B3O2F
hkRuUIx+cuY52rs+9JT1uDZB0k/P4US+04E3wUPjEEkRxUYqsWW7ZigY96R4U1gJ
1cSS/kqDUssmfpJ1s4PtxzrN6WZxVzk2nI/QqYeYya33EB8LH9un2aYyp+XvXPWx
P0LcAqTv/RcVRFf6gKCX3g91+c9yXBWf/SDvUHjtiMVcSJao3ScZA4hfF5KQOQFj
qKY0wvMgSK4tlc8ejmCPZ1h5SEmx/qwRWRaPNYYTuRIdEEVwULG2mi7lS/g5SWIb
XT6QFnuGwQ8BF2oepJkQYr51yPmjL1f2LljpkUnwuCoblFZ5kQTei1R6B/WrmFmQ
Bpfcf25w/Ez3m2/GMVtGqALv5YrG3szKSnD7js5p1yzp4dFVH8TxQR6kOSncGdre
+EMdJ/oaqZLfgnRRiAMVjAJWxGhcc8wEOXWfRvvjdxovEfAuRG+UwBEs+JIoYDBt
81CxWBHmyetFaxTaOvuHtbVdDdQC4AJndP0Tg4bz/1qMc7wZV1ehdldTQDjbjw+k
3LKqkAKRkgxSHsa6ofO/Laf7neLg5HGeFXqvdscSJmmpSxo1hFu/ewAA13SxMEn7
rfQUKXHyiYYrdKvu4VSOaw6pVAlDrc804MmyrZOE+QtuD+tep+N1w4KedOy0ANjS
iMgLQm2utPaZcV8YALvkEXUMTQPnaQBFfjqebDM/ERNC4bokoMrR10WOMe2fJJlj
w7ev62ok7zQ+ll3GKftfHI1VzZgDmrcnrTKKxqsyX1PP/2PigD2GnNSTB+nIEEJl
NPzSwko3uzpbDlPZ6GoIiR/ZYKzvDYburvsmIhwIXbsP/9yJEozdRb6uxqr6lOwd
gnZLAl3M6ZA9kmJSzYqFsQs1LOYmH06AHeIdoShf2Gj3H/Mk8+odN58Q8dZ9rRG7
N3jqF+e7YB4vudAdpn5QtynSeWxR4npWOkAsGYGUSokxz0TMiVHbS79pMzfa2JxL
PuWxrSEAk5pOmLnnuXqGCnpySopJO4+baUz9HTgrsifig01S5boQqv5HnulPui1L
SdPTgAyVFnmTjRJSyEAniBmc3w5kEKiin1Ayq6RrKf1hnPt+fO3moNiRFWKmhKTp
5UQ7xzU24RrBqmn8waf/wDqMZYEyhWAYOTYB4K8EMNBJ3Ss/GXDJD0pGOLQhExss
aUIkI/vDHLfvRep8hafpFldPiD8aHEX0Vh7qP1fKggyO65Nzx3aSL0pB4r26hwkp
mo1yEqlZ4I+s+edGUFi7QprKbB1b93sHVxfGblacSZ/nwRDFo1/1jEEj1CWSGVVK
bDSnVeSbUk3h3kXcgSk7jwKQqng5igNstHI6HCr8q1XqLiTYmcsfYCP+2tDm9QRs
lSKE1czljVm/Ndr2t6yYS3Gsogt+TNTGCBLS2pnRposMwxDmYhbM2ZKBd5Ua48/H
vMUcjtTYSDtMXwdOsunuDkRTipETgxBx7iUsmX7rm+hokl0BpSsUlwDNl1hXVxVu
Gxm1cqVueLmrFPwKSdKwJTp9DPYPPrvmXgMdEFwc5aUp7EPBsqD/lPRchtzNHK09
UGtUoCI0l/VgKZr/BvEHzc198olXMZ18kLYgMXPL6QFw4NZPGWXBl+lGVP3fHBX5
rK/qK1oMb5YKnOHUB8AcLCpYP76adMxNnao1Sf+WKtIGUUWfZ98b0muGC4vZ4xAJ
tpsX8h3jm6nAaFk0ahDcqkbGy70D0TKX+WdFqchrZ+fokPc+ZPhlP/1ueu3IvmP1
4W6QZcqMZsmKWijPNWNPc1Ka2a3PhMxtS+EvJsBYHJebEQAXzZkXi4f2cNBrHH3S
uAv7f3qZS1SpCHgPPpdzGKxJy+x/NXQt4FzDKFeHVtRfaBYl2NuBtV3tbUAzkjyH
MXwHKUUfg115voB8fI78pRTTiC7dpSzp9M6VGqrtJpqwMqjDu7Xh5/WGrNKitf08
G5pyXSMGN7AigjvMY+l4GPiIcfwbS5w/ZEzk5h0fN4m/MRbsp399ei63Uqu1k9D6
I3QvoHhABWYvT1esbyDX65Xuk+Q0h4KBz36EKbFFp6mYcUw3fsp3VIhjrC5hKz+i
tvupg5lHAK7cdY1+Daquo87sjTVmImHPYclkD7JOhvC0jjDpXWXFEipYqM0aQAGB
P2JFkk9LmtzeXtS4blFlG9Q2+KbLB7ne6BJVR36f73faBG7S8G0PI9tQGPPfyT/s
O1msqr53ZIJhdvQYk6evNx5yfNOZF8zDy0SL9sauY/JgRFbflGcXYZxdIK/laO2A
sIwzgRMSW5dz6ndb21uYsp582UFo339CV6Sk/Ns94kv4E/OWf7mHFmgPrlHgXoqI
pVBvzLwzcRDa79Y/h9z8hs2JtswOghhaicaGAGsXvNu4BUstqqAUg9u/KhFZFDbT
keu7djQk01boL3C4J4MoOQ/w/gO3pfPG03TQ4xIMRPYPduNqizXhYFPfwBf8ODtt
rzr4lPGaE6UgbxUWEXE5RyP3iUUQdiwTwp5H8tjacjKLU+5VX2eurWm1wk493cv8
Y3JBR6cv73urDkwMM+MIz7jy4RIU9F2ngpHuovvEmgzHTosFPFyC/WaTI9vT0lj/
yCA3djjSLn4SVEXVUX4TKr1Mz0TOJrZBZlQH3aPOPY3KEsMCa4mBvQ7NrYNvM/EJ
k6LUsQizV0CFlwzByBr5mIZlBikTEa9SCvy1B4FldU7d5z2PDYP/ful+26e9c7Rg
7p/jri5GDxnGHNqapwTGWffTjU4AT0PvDJlm7RonZmMrIT/htm6dwBhPfzL6Tiqt
uX+eeW8I0xKGcibdREcBzFezIH6IQBE3Q38qBiqeMbXU0jiLzR2VUsow9albbi6g
Sy87cJz2U1VfyqzJ00GkpQgDIxSWBjgCvz7iLwLhOCZkB3QsG/m0mDDyW+L6aQXk
wr4LRFV/Ejm9/hzALHBew/GKX+KI6P3ZJi7qipxSKrKWazpmwxaUBtMN3S4wCml9
yIBMPYEbYx3ZYnEjY1SdW9Oy5LnsNp6zBA7fIK6GPw9JQ+KZgN6gx/SodOxzX4Cr
w5eG1YN3yp5fXFb8MGyQ4zC3Q4994WacPuRVQsgCenxT+SRQjjhw2bnipJ1Cb14Y
3y5QDtqJkEtoQ7+HQJjwnRP6oc1QIxOP0mOe6t7S1Fa7oQWkhcwwu3FetgznqcCy
FefSVjtZUPf+85vXSnjuetZPFHFb+9d02n9bbQ0x1zCyeInbJ6EhVrRuF4xsq56L
HHT9iuRTVKmrgp1eGQl/22Ghn2A205dj0sgcUQD2uGsXwc1sFFDxDcdVAUA1Vr3z
RkNTRyBLFnFtikjOsaUoEWxcuXQIi0o5vxUgCsPulB9AJRlr2K4dWbMZsp88PoeT
Co6C8a0GAv4hjoJwEr70YmS5HAWDsDXAvO/cTJG6QX+KKzVrUqeLTkreKVzawN1f
0o+rlb6Cruu/DdB4ZOhNkhcKdN1ZZkblw3Vy0iGm3BEZk34Nt7ZNfdqPPajPKJLA
5fpgSuDw5UqvPaZWoIb5M7cviFdihN3a6QQACGZEc5T3+6sovHvm4mMdeXDBCP/s
024grer9diAEougf4vhEVSRLpR9PC0XNDazbH6zMKVb3xNrS4xwxXVXrflJyIdk2
Ue7iqMEAatFGgK+z5eAg2iMn3//jP7Gqdk1lsBV+FF/srXNPMHc6uzScj5kvfEq+
AmKlQu+hQRykOo//FRF3eNV6HlcEyZ8AQVp2V8AtGIpnJIBSZtzCjicagtDflwPR
lc/tK7GNhpEeUqDcOsBxvFYhogEk4JjsUIP0IiQr0+6C1bfjL+ThWpZn/Wz/6Uwa
zsNv5Ly257nJ3qs2bo+fKWDxsSwLfWnDJi0s0qwYBv+65mghK17GA8bmlTBJDW50
ij4c+joJrOTrWVQkyhUBKCpXbXovJITJyjYNUFX/gTEFP01SG2YD1fbNBP7EWDmv
4f0YxCY9Jyq6bDQ39uch2bxqrQkEOckOvcOPqaVIPRpuJGWLmwPqroQgdQElSYop
ame17IpVs6Fvt+3EQZOEO6Gdm2ZKWumae3Yi3Iak9VK8zWInvbhW44dqd+VaOEu4
iyYStib9R9AAXh+8EZzXNNZyg7wsQdp2KBLnxj+us/CWOXpf32Hf6iUmUVk/URmz
ViLLjQyq+kwlkbhs/962Cr99F0Lx4wFhf9LD+0QTCzgixS0Fng7NpfPLI76hkhQn
QKrJOKuayj1czniGzrlyPbErOx12zQDpnDLpp5IqiZC2sPRQ9aRAkyAFgPdnnE9K
VtrP4ySd733RgGnMXgXCdZdEjrGeFT+rdPTgyonifDGS1LGrd7rgniVcFynaS9np
m5Jh3dzY9MXa6cZfdo3+vZTyYkH8Iaq69RIT6ER8g0yq8/qZemzU5/hGqwdHdV9d
aH2q90viC5hxuqKK+mtEB0IvH6U6TEspSdYt+NzhqNB+ys4FNM7D4NMGltFKVIjm
cOxOsz1+fZWzE9UxC8lJ1nFxGWAuH+MBVGUTrh4lPeNy7+HJKh1KZvM50f4IgqjI
09ILA1ldlHTdjV4EFeW2hfLPZEqa0MSzazX05dmIYFLH04E65hCw3lanBOFPBVd6
lgDaqeacw/D5oEsst9iMg9yu7UGhpfcx8VyegzKI95GBHuJLvuBWm7jj56aZl74X
p0xux+Az9DUcx3a+g1dWTH1m0mTx9bLrgKB01oN/abZl2Ajojzi77JKZ5cUW1GGh
lOY3JGjvCaY62gpZ2mOT9LiWqXH+1hnf1iu7fF4zgdXFuHkSHedt60iVHSJlms5x
/hW8GgSFuLeoQxsTHCPtiiWOGd0YRHqb6QjlomAamPADcVn8aYIua0flNcxZhcmQ
i8l0cicN0qqeLMNN2918MlwwmwwtTEw4wNjY3PFJwWWW+aLXKpVyXJ1iBWARbBoQ
YahzWIX1+miuNwvyT0F7l6rhygtTh2Zjt/B3zeEQBvlTlV9M5RoTWEnuLD1fwrl1
z2lUfgxV2Pcxjy+g+vFaLDHkPw9I2uG8FZLbKdfIkCudeaU64dnEKvSP7eKVP0Eq
EdV3E217vVyBro7VeVfnEzp5zbUyuThHV+pmbgzWssodkaOdnPwho7I2oA7ZY9zM
ETuitKG4LjZ9NTIS/B1Bu+oqglS9upFyVPwPU6jGhi4Dfh5scphLxXyK9amtrC+p
3MraHv2zeensR3C5K/xkikXAyeG55pFsJcI9IWEMovbSu8g8Mv2zS6sSoEqaykci
mRoaydTs1Qlwx0jeNp+1dONoUBLOOHtqg/fik0JirNFs6DTBtJTYALw+Z5q6cKPE
GjxL5dV6ZLkb61oVxlYG2NS08J8wC/uoVQxk/ugeL77Ema07hKcdGgSqxLJGsEWY
kmYvyBZhskTN45fpcPooS6PgiLHzUmXFJqxI3ltobae6hyIWpnpgXBLpQyDlNfB+
1U/mNEZ54rf2az3JK/w8DhYBIxqYahQxs9ovhg70VZZtJnP/5Qt52ESxB53KW6N7
BQ7EbwNvpyVrMOP+hVUjR4u+uY4PBu9FcX5n8XK34LiyaCs+IT5lWKCZc2+M6rWQ
uU7pn/0UpKpbDuAIuSLmr+cVPgoF/Wx1LKMQ6QA81CHG0zscnavWEpjlHnZ2SoQb
WVPpMMewqMZDz961HbQ9A6csP43GZk02kCquZwut5diLyIrp5NQeWE4wZYLcSGtm
E9AaLnFr7Z/GTF9Ce0lVfeDQjBQRijtOY/OkCVKGFYsuEkPbfglFSIGaG4/tauQJ
AMKtfWJ/m6OmGHpHPegU3ORrLnGKzZ4iI7Zl/F7tSIs9PMvtVHJPKevehF/Up38A
PbDa6LYtMKxLeFS1ruDIn9BJuCnz8BoLnMVHB53iHICh5SHEx+X5xEBhgflBG3Hv
FoilN2f8LcO/8ZUHRC4vKVEL/OQjTwhnmx1iK6Q+fpcvGP6W+9I8rTAHTAIFnY+H
nDG0ascA4QF5sssEUM9jdPzn5h5/9zrjaWSFJE/sf9VYWCjX2atlVsFFygUpVzcp
1SYspXBXOsQumiYpsPLvAXgNE6lSNekjFHKz5Lapn3vXJHmojMeqFY/YBzUxflzL
T5irgwh78kvAQuh6oPrnjxuDrokuSnCYZ2MGdGD3mVwiLxC41jF+IryQJQ9ToLu/
ng2tMYzOaafSO1kxkD571+0hTFA0ypMuwMybw+2y/Q3ev2xuy2aF7NvaOT/zx4ue
zzKVClgPmPGTzgNXd//nuaY6sIQio/WLACfySBasY8JdFhKz1oR+ZQ2p3MbkDPQR
dS5A0NQqIToo5g2BFO69YSNQM+T+yZXyHf5eTEK0s7xpbQJw3UV5BPV9Z/STfGir
Rcqm3HePDMJq/tAuW6tkb631k8RHhsZEXFT01CuWO1FnBUKmCtDg9mRAlSOn9hGY
XbhGdKIyIDEPLnMLSY2SheDYbfLxytUU6nStApOSfY4tvSg5qCwbHLUt8UgMsBAm
zcysyB9KSxK6q71sxxewddJCox6kRTCTIa3yZsfpTlzf07YYZSWMxFhW0f0m4GZu
aOHuL/Jb8NYS/P+lu6xG8dygKQPTwFunjCTBxrbusdZs6UvL10wfJFTktuEfmZVS
MLtaG4Hl4i0vMaIsJySJJeQ5j4NeWbD0VL3FfPtgDbXq54b4O7b+AYAWdIGNIPAh
NaZihdrfqriG8n3iS/0sJwLqVHJ+9RDxeJ0E/iTSeS56vyydIa/A96M172xHzpO5
JddBGWciLLpTEI0A/shiDrzMerPAzR0nldsXt2S77ZhpSHZDpiIAvTU7zrKYHjNR
4Z/MEu2gWxwLKKXt1qrbdX/2G0kbu6IW/+8J3UaZSjQjB7zOIFS5zRx7N7xl4fP2
PWmgU1Sf3wefYHFLRaIJ3olXc7vCiBwgnjDWy+74fw4Jy25SYF8ZMMi3HWUFDvcy
coJNYaWlMS2lDZHxe+TzQ96Okco1F+Y1VHHX6xlYOjoBn2N0GNx294nyGfidaRj/
5i812QneIMDmMSSNZO45pwdJU3awfUVMAx65Wp5W+ylikThB2FfDG+zLcmrtxApF
UPlY9g5h6+c7kidASYaoCfsZb6rtqW+9JcUhpKeGUxyjVy+BIt/jmDT2cX/T/rdU
NzivQuWEkMvt0F/p/m3XWASkmsdXAUGsvT7qgUlE9fXt+g0DiV13qOYbKQzUmfzk
tdeVHXgHUi9lI7knf8DYKYZ6iy0iFCT8hV/uvcw5/9e36GlDgXFyuZ/9dnj5raLD
yV2TDj8gc28vghLOWz1UbJs9FHthbpiXFfrSoUit32iR07ot80Gi1hfqZGGnwFQt
X0BqZYxfgPqn6irScKiGu5g6tiH3Mp0N0PbBEKDRIzy/RDz8E4Vj9ksVAbFKl9zA
fL8FeLakQEZXPNO0xD0uv5lCqRhvEPRxQCo4J1Il15sQoctB0lKkzsmLQJUUvjUT
2ufgylEaeJ7ZhuFXVKEoFjvoQ7PhQrVEfsL2rJ/We1dK1Y7Bg/EOYTXX5dqkvlbk
pE6tH06d8J9U9B1n8ZTsrvvvT2TEAVyk04vWtoIs02sTqNd0qZK0zQp9TlGI71cI
CBZGSeUu2f+z10aKzWw0nz8BX/fEGR4El8NwqTmkT7Bo2GYPLE/eNmHX+TLAI3MY
FP8usbAqyhQE3FMKotJDRGR2TdjEYxp2eLo+lO4Bbo+rMg/E5Fy8Szgh8ADOV8kI
Mjc42B5GDbGkMrAG+ToIF9mPozNC0gUcGDXrZgj1CgOxNCE6ek3aC71bK4MR1oCU
4/LY5wFn+uJruqd0UGWx4Dgs8UIxqAAJQ4K8mPdYZa7Udow/nsBtL699tBJ0ENln
rdIQgqnaDArT2cHML/GAP+YH8NuDmUy4il345aNZLoFCoGFJ7svUY8ejIJLSEVvf
fO+bXzIIyG/xDj/oyuvQF/uzk+g3TaYc3Ko2IvQ4jS3XQB1XILfmcvBH9UC5Lfz1
JM0isCOzRPdYIPOhSMg4GTNt2/FE+jc8P6SQp6jk4q9I28rbiMuRSA9D894KD7c6
E6zBPR1k3op2igy+HJyATxxmUwaKiMoIZCgLk/wmgjsg56Wq99HKz9I/cF43peHB
jynFeq7HnGnbLhM7RUG4zV/bTlLsoUuhQk+FpHJUvQfNCr8oWLlYCcNaUqOIMNQI
xA7iktFel6I4eMQ+jP4YX6b6h7FiwqIanN56Qwa6zc3+GSwCE7huwe3H4ZvLkEpw
9yA4CjQNn2nP4I2S9wISn+7FZ3RhWn03Lr+OrGrwlFYLIgJCOx84tJUFYn5Ho4uk
kphMFFN4vzB9E5wCTViilfaMuXSf2XE5f80j931SinMRJBPeA/xHDmwfYv46EUs+
qeOoPCJ0FgSWaLnfKMnOI80tYa1jfnkoTOmVF0AuVS4JIrcEw6lxWuab6LzB5I6i
A6A+qXeogvxeqzOdLWSd42l8bT3XYGZSgwOaKWn/bpX9WRbmfXCCy/7ncKPBIULk
dJmI5YmiZxZ1+K1RQJgQzP1Kt50ClG6vw/qs8XSrkOVyPAz443W89GH2ryM5+UJX
2SKS1KWEzc54RSR/Z3YJLzcSe4W2tXoi9tZ7ZmoLZaJaijbRUQuvqxgckBY+Eab1
NrKnVj8ufOxsLrbZyZE3PL9IRJIG9Rf6Jc9DP1g9p6JsthODHp3joLTnr/Xq2jco
syItuTZm5C+QlCqHp6eXuiY88gmOAjczH4y8bJle/JI1nyQzrMUMVcaUI7Wc9WPq
7FQbiIj+gy7lhcqk+TiFiLKrvcdt+c6WxeEb2C6ZIP+IBV30DPfNeZp49ymRLuZp
CeiylTK+FhAGFzAI0Wqg1INlpsdoeRKs9iBb/jI+oDX+pgFKvRPDZp2ed+mQi2+r
xSHbuJ8TgB+ej7WLT/S9EJPT3ZLwaJ+cHk8CsSODVJBm34L7LZY4DFRepj+sSYaR
LQlikwaLLKinHRW2WD8o3Lkqxjdn4UghEuGxNmrX5NOXT55WDaojhL19LePc5NHZ
aD8Y1G14yPNs+Rv8L+etuUC3vwHeqYGlm4+qIRW3018nkRT/LEaX6XiX+DOSSA9M
U2K/9H2r2vtgO3WA9S4nGyHwwPjTeZHkSL3RGciipNAiyyp2hViPrV6lWVBerUZI
xu+klceNk6eG/7gpT1R7Nx1pJmQIqo0JRZpk+Vu8VyshoLmFodzrYAFYSPd2qu5u
wQVi/NtmxuNh8O8jsW/gW9G3ptwMz/Sbfyk60EYN0xUS7uWY5PK6f3Aa8DL4fqTZ
ulc5y0cefuj3fuypLVeNjNkLGv/MpLLrBmAN2rsLJzUcVAav/pchfp9HKKxeppWl
LEzrpnKmxSF4yf0Kb0uKxccUrXkC87zv9xxMCGgPM8OcK4HIhmcAFrBLGIJBVYco
780ECKS+QyivQzQtChE499LfrZnN9VOj1Jy0d/jFf5J+5J3OSCSLSAfto5vq3uzB
PZf/tusfi6P5rApr+e3UbwSq7ar7nqT9xtB1S275GQl0HrGXjQsls/F0I8vJ11NL
h7mQFxj8sVeL5mz2WBKxwL/HqPgONKg+wpdWs1R099Z12Qoub4uUGIvPA95KmenZ
VizaOKKHKGto6cGAGhyJJ88irU1bf7ugpqln72xWeXFx5mP2h8XJf8OZV8gBMo/b
6MRE8c3FOq/7QYxtZhcwpAXWthOlUyZduqcf+Pr6vt3h+FCTOcAw5I6MrKyDsq9X
C3JPQKilbwK/tW1cAsDulMoLvhcmjSV8yhCliQVuSqCHeO/SeQBY9pfmJAtU59uE
QhltdHXWrWWNJEYeiZwchdkG/FKkGv/f0cG81MENkAhR20AXfM0DXum37h6//Y4y
BUcuxO+gRRNPtHPrDjxkXT/3/EIJ6gICpS0jTmk3iB8wAygYiFqGxB3SEcqqW0OO
CyVd5RU8THCbA561MZsgTTGfuuswJe3CW7I+c9RQseO14cduHGU9umFeqLXyj2D+
afNCeFTa4xInxu68yQkuwrE4TcRlYqHN0mT525t4Hougffi2ZhGEFPulMdGsseMv
QD4ltBhdSFKVZnmVUrYGMS0tLu+yJKm596qoqxfYqq/HQ2qQbQK+jmygF41w+fPC
PWVZMY9qgRZWBBn6xUItKZyR2tqNGRSmq8npyJId7HkLC9fGDbSrM/ELBsf2+B4f
dWEtpsr9GeoIA/q7S6/TS+Cs5DNp8O+5YdUTI17Zd7m4zI4k0r9zsza79PtJOAbO
bQaaC2lT/i7WQRTWVEytVzDJ2Sffkul6u9dvJvxZLLcPz8iVMUfgSraQP6cO/8s2
Y6rIbHB/1RGlGwcw5vq9GCbAbvNlPJNwZIz72wFEYrZx7L5Z9lwCDWaSd2SMOPoZ
1ORcx7cTc+7u7ooaAwnmS9MGXkBrFfWzZtWCTRedf2LityCsDe5J/TTc+EtHWkq3
zpjmafr/FuPnGNzepzDdSsUkck5YydIFIlQK3LWKu/V/VQ2GsxXLG1A8F/drkPIr
IQsR49Vys30VjZnon8yApfxpx6s/kdQamgILo58ph8LoIkreqyyx467Llom09MG0
T6fJwzo4OdNDlNy+ngav0mdTve2/MCj+zXYh78l31oJAUu9S1Td7KFrpPIcTH7ik
hN1/zlbBCkZKFATK/cHWUYEWCZAtLlcuQqLcbxLSfXwRbOGNu1EvHNFuy026lPCy
rLZVKPJqbl2BIjsb+++q09NwTRfWINeN3hJIulaSzzA5ewPl6Hu1HVqczxdI3blc
8QtlzAXGlemnmRKROoMFw+DfnOLCQXVi3z8ooPAp/wB4KQNdPdco6lY+lhBeudbj
pX0VDRKkU0zvN69iw0o7B3aN1wz0Ityl6Cbpx1eFOpRN7cmi5c8zLhGgloR3KLvt
YovvrHXcZ0EEzjMhjIf94B+t1L6U7BvYLNlMJbHychtHnAvArXtW0ghaGdd/yCQT
4j3k/td/+rVppqmjZvqCFa7oHa51EDHcArp5ARCL92V9SLHGte8xRaZZVdJl83Y5
/oaLnHKHVhUfzU7u+w4MECBw2H++nREGWjUjZf9Ipr2keT9VavF48DsuJu3jIbYo
ZzJCnI2Aidg0JFG0IP285PMZVpvlnPXoGCcKDGLcxP4u8CfcNj6QSmuJUZvCkXeI
5Zs1g1ixIHJSj6EA6+tdY5iR1ghIHOQKYWI3cXqf44VX1/qSHdVi/w/ThVgFkVfv
zzl+byFoXXqO5M0K5jWT1QPfWBG/46plYyEFhKXmVio05KwjWIbO3AJCRtWWh9vT
pO7aupKfxQW+83VPMrkdy4CTOpixM8CYCEhf8WekaXO0PfEI2n59PoyQNLVdunSa
Ne+SDy1aJF3PGmIGkH57F34OZbXiH2OegxjqIrpUHEnluclWy79QHgGAElpW9tSL
xvoJDIbprE4aJK1UdMbnCrlwEGUE1clDjnZA0i3edjypsoCA6jCCDTfK4D7hdEZm
NxknE9nSEdvk3kg7FekgM8z2tZnrRGfISNQHVrC8sv9/qam5kJtVxmcoaFxzzOXb
HxhweUGPR95E/rnXK+St80BOjGMt93dUwgQASeT5j4J1XiH5b2yeH0fIPTKrgn9M
fdrDmv3FKSfzYOcmzpIwFiEmfvqOgx88izmW4CJA9gDTnvAubBVi+eqTOwPSQNB1
XlokROl8whLC6rkNfB8DdChwNsAa8BeMbH3hi+iM/S08bQUrahXf4jvFvPMj4nAj
RDobpzjjv+WQwh9zbVt7RnjK8wVhbvRIbZF/8z7cKnNS1vDsCBx9SPjDPAzQ/s6H
tnR3kzsHKlLETeDdZdsztG2/pPNYsq4lEu/wtbcWLT4lQIfTzSFZd5PBPrmk+B3A
0bBPZI3mV3JUJIwETsyjW5MEjjo+r7C/dFE54eZdS3rhrLn50bL4AudWxJLj/QVE
NQ8YkNrZDNr2T63Jbocbwi2snWwQXAZuPRmK5B29CxdCaxBXsqQ9U9WvKotc37es
87dfJuc79V2Jd/jFgnqPdXhe+tasqXX+eLbHwEQa0Bb1/EYDZDckDT4Ss/RGjcpH
iAUIW2eQCrfHQ+4kFnmKRfGiVwN5ftNGG1fHT83tNZ8tS0AkipsbXxOvusoby6sU
/rUQ1/Dv32d/J90Kwfic+tIc5el9D3kiFVNHJuGRxplTb8WamG86iAD2UHT+WsVU
TTCRkQ0SHr2yn+6m+rJIjJKXsQKW0gMW2vMuK+09fmsUEQrnZ16QYUdMtmnMt1rH
xagdSqH2eGhAGO6QJWxxwjL6lZgBFfS9psO3rp3nChGjsw/pg49FwLyuEVn0mtD/
PHp0f0dNhq9vY2y+gObKJKqEdruARyeP3A3H1Yj68UWQKN7ylE7chAKSF1pG4ptI
BdhYO7mfIldm96b6oVcymKPy1+x/6HuYtzMCYQdxpi76D4OlHa32EDju8rPhbWAi
uqnVrcpTsTJNQbRG5cL/ZayfAwJL7V5TjvJZHtRoSHja8WnNhAPA3u+yoa1MKpJ1
HghKYKutwHJlV7w1GvNurmpKjCMABhYGPYSQsgXhifpEwlavz/vJo7F/rMq8JApJ
VeyyfwpQ76BzT81XcrVal6tGSoJGAWd9Un8ZPV8JLpiEjGjy/C3839f8C5aAWxyt
axnogIb3Uw2ngZLwf5pKiHRGsct8UTGJWaAXBvh7/e/NyEt3fupGIueUS1pcBOWX
tOmpiCze5uKKiSMSWT+8j3Z7nF9ngicPRY9MdnypUkLrC0ZPkS75RzriLWUr7QB3
QcEA1u++XhwQH9sup+kr4VN0shXsWYxDal2uyjRWfRcNmCJiL7X9pn4LcV4AfOnf
OkO9fHtB3SbIdQ1QW/ZPOvXQCFOsraRCGR+5VkP7MlOWIGR+prtXZJmoaZAu6Nku
NwA5JHVeZUlOWx3L1xVyqDWpDVEfv9vdDNRy9e9mq3eibwT2Sgc2gtJGOqKyu71x
XAS4xna0+xhfLqHNEWIP6rjigv9rTIQ3darjwGSi/AOEEsFyzSR4t815VgzzmfZP
BUmzY812PKe14kq4HkmZxryF1iAo1jDh4w2Aczowp2i7ZdNzh3n+xMGEBagA8VVf
yJ6YjF74JJRtz7yMwyR14lT94kIkosnNsMgtrHgQTZeCdtc3YaNZx+/LjR/7dChA
u3H0YZ/vFFNFn0Jb82TUlJbirLulW7I0bMkDQO+/+opU4Hwpg55Exn2zlBtp8KBC
Wj+KSjYqkNmbtFEh5hrZdaS7a+obrcBUu+jKfGB9Nfqc3n7f/2fAJxw+Fw9aGmBE
Xo1Xj6ZrvCONhNzd8qpJ74gvMcTwiAIUHdWHJjAuUjAORikhS9tzanp5i6okciVT
dcMryDoPNqjwgn96hct8SBORyscgdQQSfR//+CON9X4u1QE4lnS3HecUyF19YCbb
g0lDmIcQcwqly23IIG9Wy3unelBa68/sfS+lJTIw0atLgG4jUAbX/dHZ06RFrZmj
FViMIhMHjdIglJPZ/idbajdikH3+Bt+nfH7RajyB6BLTrW95yN8j3us0U7iOi9BJ
pL2InDp0KORlNOi6uyduZcx09topWUxNVtEczvHeQXkk/Blb6+KnWEGMfIQZflW6
l50//Xvf0xI1bhSeGOKE2f7S8gAMeUotqfJXqtBve34AM57Q8zvVpSBPyPyupg+f
rUjwTb7lf8GRW0ml0uK7+0JUv/2Q9kQqsh4eHZfzxqnQ/qD7I4MhfdHHNYPGFFE5
jxsgxNJCHGshWXTmIFlox3q+JZUYCSfHBeEDnN7/dAmWpGTW3FQFzrezgT9FXEjC
+NK73jzqZQWepLbY8GhMuiBaSrP37HbZfYv2JyPruKM51CZC9Ggll8B7BZhQLYEp
EYVXstiSNsX+brMUuMS+XeK3Wd5VdPwE+EqGJUlBS56L2/MuaE0cZdHxJrwQKRAA
gROlTgC1kUBhcYEj+YcNXIjNBKr51jPpTjEzC4eQd6pda2H1Gw+6kZqU/rucLtxe
ePj9U+8rmVwT5y4VE1HNned/+4q8DYRmLFAk+o5YLr5E8IZ24xHF3zDZVjxOLnlJ
DhCnB+xqnV0BS4eN4hZIsMfOBMb4mhrfmVFSzygESqzu6DKT0D2IhIdbLJN/HzIj
OqGiKyXL2bG3594tyzWZ47QxX7xRUjSTjFqpSxAt3sxnTmgd9WkzyntSEUNieA8d
w7OfU5lE+9ATZUvWMXRkD0Ss/LZ4Is4GNQ1ohoCOuHNLVLPMup90VG3fas7/mXu4
Nm7j40ktEK1EhQj/+blnggzWlGMyRc61lN4yh48HyAItsi0Oobdd8ZfCVSipYbO3
YdEiiHmES4+naN/IhK7bsM3/WpULXJ4wdZD4nfs71etrSGTbmmmjmiug1xPhTYnw
INF7lhSqBi6EtWSswBZ6w9QpZXpBYezW5tYukfdCtTdF2spk3ITFl0/OiMT/tbGQ
4UOBFVcK6EabqwD399BTOVwrcaO9MBGxAyvtdKhXx+0F2qMdcsv97NFostkvW5oK
auvRcFJyhRPoihEEdLLBj7JtalFcbMEhJgmM5DAh8tr7QXI72scYt2tB7Uh0nnsJ
lOhztNDRe0Gc+QzgxFsCc8ULfXqJNCCI9m8RU8EWVfThHcbczuEOGo1P9exV7gYD
l8RxCpTBoWFBPzBNp8EFk2ly+2oaLorg9/rnXGkTEAXCyl4aeeT5hSMQCwYYtPfi
CtXmMoRMhqiWnWUsfgm1f664lAClipacyRIe6DpCCXhzNFk2ZXPGKJez88ZgEd5t
YbjAQacG+IvjT0BLa8pdvKr2272s0BmiewFnttIkPn+1ckixsv+E1XQk4X1cXspQ
7kUfm0Y7jBRAUO+LpVt9kCnBnqvCh3gas0tJgSsrUf/dWt/UBCpvM+PVVwcoXXQD
A6wEgzFdAEoO8EXLu3KvsVHtWul8Sg9DZSOATBGk3cwFn3tr4b+lxa4QiE39Bzb0
4XmxpxTY+22tdYicQRZ4YVt5jHbwy2GS9OGQMzvY+NKQPGjmqmD2dVloTq6c24CH
iJg5NebQLHWWb4FYFLS+urnHYVqKql1PGPi+FFaQ308/Xy7Vf2lR88NLmbW7bnT5
Vji0q7iqm71Ef638FwZD61j5BfWCZYAkA7zeYv7EGjFUw0/Qg34LdUg0Bf6BiJMp
IpVWeVJpxKqt0R27ZNokv51RLS4TO8jcaeJyPaZTWmXeDAzr0IQDf4x6ump+Bkkz
+UAPMc5RV+GdMfVPAi9srNU+BybO6nIXYOUBzyXGjxrCHcOrQfHLyqeFH42T7a7T
vOb9zCvG+XrXDf1hcTNc1GcUGewkl1uMCGColp1q1qtmxdrUPxcHO5dUmV4ZK1SD
gcYnQ2uuArYfS1zafA2IqR7hWpPI1zR/RgHCJK5FqUHbrWz5s7R82fZWpRIG652p
ltwv4wfC6BweLuyZrYrCsxLfmguweq933Z29Wze7WdK0JJe3TnV60Z7pKRhEdPMY
EnIg7+JtVCYkqg9n+TwdvjFZFkuVyz8Yd52n6c6MkaLtZnSGsMtD8Rma+82Un8zq
cz3Lx0I2N4M6VULReA4pgBNuaVd6dlHcNX095wPucr9n4rkPp3pDEIFWhf8jKnxh
JYzYaj2tEk5gH1MaurWtAS6FF07EyeZkCZH1L6xh+3t9yYK5ZboM6aJjOL+8l9xD
+ARP7ib1/Ef7EH+JQH48gWzd4HQwpWIr0S9o545N1j9QbaI30UJQOzVLukyfaIvy
G1sVsCetPFBY7XlJ250VT0uzx0vU1LwsPxdt2LlXUZSZMinTSsmkG0XaI1JJfePz
5XvfLGrztlN82fbwaXd0enJpME0bNBI//w6apWMMGsglSpQdGklXbvpldQKPEomJ
hHJxpn9aKJxWVQxLNYi+GEjKrjYDYOUeiHe1MgFxA3tRqgn529jdt8zVYPUGAEL3
C2hjxpx5SKg+4QpvucELRIPrr/NkTEVx54e8D0rE7luUcsPkjKHwpWzVdduTb0Tw
6+bg+dKOZ1XQGnzB2QpcI6jML4k4v6OYf3RM0StxVTAT/2oBkvBDZ3yNCrZ7X3+K
vKx4KXFMVAXrDhcucE7TgCNUuQ4K2nXbM6lHIj16Li1YQ1kGmt71uc1WyAZdiXA+
hLzABZ9np2KbHxaJMiPhOhJSpcT35xmK2Z5GAqIIvijb3368WAgnRTWqG71Y7z09
gh1CRV5upyOQjBmPgNpnqsQBOMq1mG1axNYIddmvZRRGLA8278ezKFtowxp2C9UQ
aoe38YXMyRPubEw1RVjlYUTlz3xlOiG+N+RILIOFfzs+2i/vitwlSdJuOMVBwT9S
OAFOGK5mzRSmGn0SaRzJ+0lXWVpuDiskTxt9B1Bm2k41FbBUb63v300GZR/XF4zo
cWICX9MuMocffQfr06mx3KD0rlFbugybFH+d2VEY+2qPdF1qQ1s8lVOo4JGRBjkz
Kru/llilYHSJ3Vd/awxtt4UzmLNyEgeLdBuxOpwkvF247oErFCXtHr/zwFNusEmq
hXrM7CCU6Dq0SuRe8ABzNNXMuVHSfBOYT+mrgE3Zk347hNJu2g5gc8MSAEF9ws/P
8kKDsN9QMcXkDk/7TqPGAoopEYFqbYdveemujXgcErzX+X2fvlmC6Q2s/Qe2xg3F
CeKhdq8EQksfpluOmdlmXgxehVAv+2zv8/xVPWpdLjUV5GGfW9h6jLN88twaokAq
ZlUlBvUnw4ttQAqiJ3Gj1VVM08E4kcjoZ8tHknIKudbrL7XxKK3L+hSmE8ybuaRz
3XKQEdkDVbp7DmuKz5UEcdxZrKm0Cvl62YZ5Y1ga6vPK7Wxe7bzjnE9B7eGzSMRU
eNboYqzVhlsttjcPKaigzylLDo5m9BfTu0TIZ5bjk6kYNggpxMFYDHF46NAfM47T
+gzIu8V79OkfVjby1WI/UMIb1hz0yZlTyOqV0W6KwX++/Ujc++I2qm8GUw5mQ/Qn
gG/JmJv92olnfuCXCwtjVnPVurUxtO9jQTM2o2R83KGseh0dL4z0tQBd9e1eN65q
y3gO+udM0OBiKhM1tu62Hi2Z75KWjIKwqV92c34zAN2yfCN85MTtWFKgl9yJSGil
Y2gxCHcB1KExb4IQke9gFWpTIRSnImu7HLFBieoMGTHpkatoQCTW+Rv0RocUP/+d
2dQKoJhA2BsepKX7EgoP8M3BsfmgvwsnEI4ImJtdrj5zfIBUDe6+SVtF9USwhp0Q
ItkbFWhVdmTjcthECcIawj8lvp9jQ3b5KEr9WzpVz/o=
`pragma protect end_protected


