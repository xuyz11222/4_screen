




module hdmi_phy_wrapper(
    input wire      I_pixel_clk,
    input wire      I_serial_clk,
    input wire      I_rst,

    input wire[9:0] I_tmds_channel_0,
    input wire[9:0] I_tmds_channel_1,
    input wire[9:0] I_tmds_channel_2,
    input wire[9:0] I_tmds_channel_clk,
    
    output wire     O_tmds_ch0_p,
    output wire     O_tmds_ch1_p,
    output wire     O_tmds_ch2_p,
    output wire     O_tmds_clk_p
);
    

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
nswCytp13CMnCDV37ezZ1KDp7LaOmafQLYqGs6LU3+rOvhGuzidaTGj9uVs0eIuK
h8H3YxEYxPhBlus5XxYxZbcz3ly/7hsDCWQBo1vFwp0owEUZfz7WQ7V5+duYfGjF
+nhD41JvZeMYElLQAI8ufgGuGkzXBFgAR/n1OAsf1VE=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 4800)
`pragma protect data_block
djlPaHJWaEFTM0lUNFA4UNV1/Ie2BhhcTp9uzrepRNwA7tvK89KfMxfp84unaIin
gC02j0OvASUjzimfUkjRP/cnlkwa7jN74oZyHwzrpOR/1mTZ82T8NvyF+/6FzI4f
rRO7Bd8hVcXSjsnkTtthLWknpPzFk5DcAjkIHd/OJ2j+SI9ftVE4XZ4FdzprBOdD
VvowvItcSjZ/PpMBxPQd77x56FCivSXNlPMc7FjsLti44NfY+NC2IjAIDdKkZJte
yzvK4jjBjRdjF4FVL6sWLtfNg1QNsTU1ODrNLw1EHzNKlEza+VfYuXaSKilAo/F5
GNu9r5UstK1kdDXhdLdCLAckv8KJA57UeCAxluHQpO5/gaKFMYpAWnwDBIdCInHW
9Si1fX5A8KU/DhAO01/PU2f6/3A+GdFUgsNQ6j76j0y/k3zIfrROsrfIihbaL+Ze
dcD4F9Rj7doHJZexSJ0DK6ZNvTr1urN5wAmBODnMTU2E3QedVb+uN/rlk7Hb+DAg
w1zhoWlg+gPc/mAy2X/RQHaboG3eqkHA3VjORaDajuWYEVWDsSBxt4XMUwO0j7lZ
Pkic0XN8HyvUiWFpUyDhkDdv9fGVJJIC1p1nUO8hNDpwrVpEzjAYLKraxeQ7Dxv4
Cv5nMaZz3NrhljtmeTyFbeFJcnPT/CO8CEKnsdzbA9aHK0HRIAjuY50Or1cVOZGq
0XXAqyck9tXRYFhL1++GWNC/syrWhoo7KQR1vEMnLpqAi0CmSk21JeFZGVLz/Xy0
re0IxP79ZqGKcxIQdnX3VsF6dSMgO8+revb8AFSjHzHwZ/GfWfOg4Ww89bvE8FC3
3QTpyFcoL3M+ajamRgrxk32Bdjci6OYsMUlHLgD8PAjM/8CZu+sHVvRriwaYHY4e
0L5CVloH22yebchJhPugyfY/HMs/Vwbsx6WJpG0C1TLjRPVdAfTEI6k0fqIie9kj
/rVclZPvwXg6Xb97xsJLTRPJcdesXRuXdUuJHEms1TIwg1PwZwRn5I6GxTxNAU1H
QIzDb/NzSZjFkwt26+60uL/VcfsVCEULzfHztRhvlKmilpIvS1R6LM19ENcXetHI
QVf0oTWHFJdoSfk02hzyR+CREejo90agY1HTCMgfj0EGZboiMwY7ZcTsRtYa5a48
ZGqO6ktQ2EpLexyayzlfXR/RMzGqRG2bIe0PUVwdfDlmWnk+WUeSn1KS6rRFlzPm
O0X4zeqncnPlSwYlxK8lF4X2UMLYB3n5gYW0GXvvV58SNo2ewHnZcYehro5PG+Qd
V4q9WzmLhm/RwxCexg5pziopWhwbr1qhh0OweURWgw0R4MkV8uxlzvU/HFu3dXnP
l0PW8P3KsD09N3EWkz5QfG9sOdsfd+vBKJ1evCCBvofwrl+YWNvkfNsYdkcpdFhj
EwnlPxgi26LRKDoAE381fYS4/F2wyTCu1w6oariRrRljPEifwQGA7ugaa1svoNd0
9dXwlB/5w59lyGyb/iwwK2aLPbcr0bCSns+KeTR+0LS8IzB7J7jcifZePOPvK0XK
yZ+TEQuKerR2tfbgm2+tJ4ZoC2CogziePOW2SfRMHoznr8RoA+AMVngkSAbonjoe
F8pPoQrlXTopTWHJM+HtFkiinIjX3hXAU+S/HXqE0HszndmjzpxDGoc3Berxoebx
xBkI+IMf5MsYZWMQulMg9VtL7Kgr7Er2NBeMotlEiHqT5WQP2rdDgBpO7mNwXPXl
ztrr3RPcjG6ZCJhm+B/ahxB2n02fxSPsvOEeNaiQbdiPsp5Fq6XcQTJD9qB3yIPl
hem+XAddFm1+RrzGHq5MIsIkmUaYyPnS+KKNSNAQCV4EZh7gCVTD1EnyX02cyCQi
cBiXDDK5ksQVkCbdBPUIVqdQqXcrWHF2RCOp/T7DZprWzPuB7zoKK1uIv02ucOXn
3RuEF9jQL8Y3+zg5jQrrqodoMLob9S/OOQe1cSNjUVK3Vk2IewSuwoDo87O0BDLz
jehjWKc4cAIEzNsqrf2D3933D9GX1nVVVCfNoonniMTRrkltM0ooaF7Re93GrTPM
P5tzLdkEs6DyctKtJpuSW7srkMy0eSXZpf8MGxTsxaH9br+zGjzygQOjuvgm/pwS
M6LYsmIFJbaUxfb01mevgvvVHnz1SjJEKG/lOVFPwSBVmxYTuWwMZdu0EeVmsLHi
9ODf7wa2gWAUXLu58mri5vvpLaz/heeZvUxAaY6GiUwZrqgoLzFCGsta1Gl97zkJ
xuRzaTgYmkIez0BOjJb0L231aVXowyfNT8XxPHSsto33piENXK2dXTtLKCdSdqtd
Olwdf6nZIAULN5U9gv7JcXeYa3zednEUcRgNaxHluvwCHbXcdLJW++PnWbQrCWxY
1+X6Gi2TITone8Ng6MVnsE20r1IWAgAhy7D+F1XfoZy0FlDwe6V13BPPUYf++oj1
ZV1YBpSR2PavXUYeAuWCrP3dxJzISqKZNnAOUZnyBI7GpIm3UCEP49YYou4Pjf99
ygpYgaEqigo63yaGwTvcM3yzTE78bHEV4tV58o4Q2cARmfzaCFyC/y1fJGNpjA3t
2QtylvFE1YibvaSPYH/8Y0KSRLJPHIH8nW9w73tWQMfLAE4zH8zdelvZSayO3ZdL
LXcVwE+0E6zDmAfmBSzulwxg4/VpX9exn6Ue8HBzlKVRPcko75Nn4T/0iEcre+5F
L2lqDohnK14ZcOIyQZ6pTJXYNw7aHjTe3KeRHzKvALfXfQhJdDItXw8DzioGnNew
FNldezvvsSVC+58ooqHwQF4yHN/6MCi0d7DyuxNzdKapk2HLkcwVVHIPKPR9IBK1
9s+jTGiqzy7u0+6wJzAkx0DlgLMLY1pgWB3cjvDcz65xKMK5iz2ZHJRW3je0K9k7
hbi2003b8V7veEF9lZMLwX1SS/t4eQFcfq7Xg9aa9R1Gl0usDGR7IluusoPNzhdk
8Z7Lkqiq9axKHcT1NWI3RHBdCm5KqG3sWOPPbFBLGUmZMRD7DouorApGXqScylv2
ohxtZ1WWCoDIiCt0hBNPfMkpAjIM8MxuZKB/neuNB0fF49HSDa2cFTQSkMraRhez
fqeVEm1QwbYKbVegpV3K43pzYF/wsWMe7X0RebiBvgomG+v/7ongS+eSbiNv6i58
CirqM1pgqeAcpPKBVogJtFqeFT8sSSVCruu+SmpiCkd8AfgHBkaqs2I+2GOWVFIm
4AH5iI+xDMQcIiyUwGBMSsoOzVt5CWbyzH/JGcsblgBfWEoB55dXjqWVHTZ9dHOi
YDmpBam2q7o26oZ+Y/jXs+OfXrBTnhHzuxQ7Z37ujx1tx4fIY1+Zh7rKeaXPttGc
dPtvEHOLx6B/6KnrmG4UyqguoyWLz+ED0eK5TzgYDlYoBN17eRwA9SjpGskbT1zd
yrpHeliFpzKWo5u1pC2l1ViPvmzW6yzF7msR6HcFTYC2KgHqVIqI/EvVxYTpFvAk
0WNipQVOuxO8t2uw49BjiOxlt/HnNXHxQGAlQnNMQV3YuIWBUKpREVFIKUjSzyAX
lfvqJFDuqUedIwrj2LsC6N2whX0hXJOiufWLcnuRWQ4APHVlkDgU6AJcz/5W11VU
YukDnZCwxqGnlAgr9dBKzbqFVvEEIhU2NExZNxLHia57BBdKQjF56Rkp130hESV+
rDIAcHVPYyqyUrIff5FK5Xa2mZ8E0ibLsnRmbbuDxFXGjMJbRYxU3C/paa/aij1J
5xnW9BfHcCufYlfvJwxRTnSbA5t7oPaX/NLeLMOpmJe0ZHsiUb+6jMIKgAKpKGko
VCoNmLN4aUkvZWJwm9W4inmsnnAMLtYfs7rDbROQhs8cG5oM1TEDWlUwUFNOPPO+
SvoY/uUts96DmhgDrJCdZwJVzcAEWSRjfoiF0sq13CG3Zs6cvu2PW+rOixQjqwzs
CC/BkRZve8gxN4C63u5xdpAP4mpM0VBPYh1kNLOL4cel74Yj7plLIjaq08F100ef
1EzDLd71n8wAn9oJyZ8DxUL5AguG8LUW73A82X37ymblMOGPEmiReyd92JRMkp5f
BYVTrEe5p+O9KfrXIf2Ypb8+KMCHtHcG3BrHQuLdNcpPAKwCLF6eAqTWWDmHW9uv
YfOLCJmeM+LDhNAzfcYHVrCLjlRNpFJv2bs1e47LpMPjbIM9pYk16PUxsZG2Nq1K
EH7+PKkIRbsMC58q0TLUU9WwxORw+rhQI/S1WHPAyNDdyn5o9/K96mVc3BD4NKlS
HfxyQn+fCQSLXHO2v6fETSwJ3WTy46hxS4DJzK3jI8OMephhO0cOAkY5kWM7+xLX
Qr19nMEbHwVzQy9jujSD0z/T3xzn7sRvWu8xFgnL+haIow2/0nDmkVZ8z8ryIU9t
wlW+6wJo+P6TVfj+2RyZu2uLI6VUWEZeyx+htI9zjgkJjGyt60IU7eEDONAXLsXO
1SIZ2hVighCIH/+ejqnPleL6ne26q0GiKw0yDetf7/qy281twCbSlqJR9ATpOHQj
IAYmmRLIWpUVRB4ObOpxBrAodJRWU9EJzjfE1rz2A7WmeI/EG4pjR7p8qxMA9FYz
j8QvToiqWuDo+MDfUNiSGixtZd17VUIHiKtnpRjceggpL60ZEvPFjoGKwC9jnb8G
GRCpkykWNB32lCG8wNhCSf5sye8D5KsAPhPPqyuCn1X8TEBhJ2LPLZ6BJej/g7Om
BDMLS/qsdYTXbCnrtu7+N5yCTlEPjZYXBDqI2oSHpTGPxbSVdk77o0QJ+bQwolVX
rByA+UnQWOxltnEFOAMT8IdAE0QPd4wCBJXm3/St4eNANOsWqLj+THNqjlQpkvA4
wQ/zZ1vvu8NEJfbOEaJaDJCL6hmYUZsippNTGq6gMnl40gegZBOihrP1DsNyZgk8
HUu9APe4fVXXKUyLKAP86jC3LBwjRwqBcb2agrxxcPCOqDAyaaRgHJja0XgrYGHZ
SKDPXLVqArFi8dfztFjvS/Kyt40qRlXOpjCdGvZyi2ycw+5hxPu+KJYNkpem16KK
rQlzHR2/K+gbQ3FS04vznoKypJhEJ5wbkN4F5HGw5DsWTsCok4CRauAw5xQv3Os1
HmBwTd3lErVB+wlBAblsnMkO1tZAeZwemYSVcsREfSKapKzSvuShrIOePicLjd2w
lQ6t+Nppq7mitKzRELz55HufQGM5i3y/r9n4WYET+vRNwbbTDOB/4YL4yWY1mvfF
vtHM7APVgO5w8iqGS+6IkrvBaxQ1a8oYmOd2qlzEK8REWs06EuP2IJFKWQnQR14Z
h5Nxu6Lwv0f000AktJCP3z8HWA5rz8nt6drL5c24rBSzoZPvzbT+VAq0wSq4/YB/
+om5TqSAECEPEKJnlGPri1pLali5IbxB4OAT43rfjNzKgXZDaubrdM9dO3EzNyK8
3QSLoEfU7uBRanIObEkYLaXU/1q6SvHCbkww9H0HzAZaa+esHqHNQGwnykZVuX8X
C28CMRhGqvRE0E0AKp2iT0mCew6q3M4TRkQnV9I1h+EGsevewihxcufry0mU05Q5
qK55fjJ7GQvHEDwKm+9NuDLbuc4HqDm9SLaj8S0JcJpD8yBIMPskK4a70L361ycv
LaURrwYSCgpjs89aPrACPqtb7zuw85T3bCvcjXU2dS9dw0FUwSp3Dp7jRC6KALVa
IZTlyzMA85miu4a/ss3sx23/OKd5dg7zrmb47ItodbJ2D8T2Fw6N9mMFBvXhzgbO
A/JluPVPRBwnSCC2orE3C9MxYLU/loxUr9a01MS/9NkT+vYy4+k3HocxWM4yy16X
TX7UTtkv1UN/XNvwYf8K9ckOSPGUEy3EPDLhfb7bjpoJh8O5U5IGV3tJYeyJ6/if
N3cZnL7MtrgDc3OAh4PmKcifUrSQ5pemEilkBGQGfjt/1IyqRx9QKVHoEsbHuLZX
vBVTIu7bXsYpA7/yxFwdC7X5H4RrdB93qYp7O6Pc1LB1z3viS+50YSRX6kvnxgEd
nyDI1B5WmaGlvAHEcmLIHoeuK/B2hraloUSfcXJSGr0IZSE6Dy3A8ScnNvjP3830
2JyruNEIaavrP2mQO4TVrrX2egfWpr/pOJLOn1z6+TgHejqHJooCf9EloR/1DDOq
RSDjTY9k4sChiX/rXuUUdrYDYR6dRRe7KJUExYp8BtuX3ZJUAYZuaeeKS4Ng53NT
fjEXklRLHPHt0wjTsL6e6MlBQo7XMavY9gs2v4CSa3SPAar1RjQoZMO+8eKPT6j8
TavMHLlrMHNFFqJ3QRNcijP8ByFHdhjrSnVmrEiE3KI1YIsSHaIU+lSao9oLu6SC
3/sxw7p5s0agAt6opltzSV1DbL35Rmx7+tM3Y+ycFuKVkZ4jBelTia9nvJZEpBeJ
ylUjUSG9wbtpT3fFUyyQClqOs9ngSV2/bNXhlI7PsxRIcdtt5DeV9Gy/7QRmOeqQ
`pragma protect end_protected


