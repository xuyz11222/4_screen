// Verilog netlist created by Tang Dynasty v5.6.60427
// Wed Oct 12 16:01:54 2022

`timescale 1ns / 1ps
module eMCU
  (
  CORE_TCK,
  CORE_TDI,
  CORE_TMS,
  INTERRUPT_i,
  POR_RST_i,
  SYS_CLK,
  TIM_CLK,
  dBusAhb_HRDATA,
  dBusAhb_HREADY_OUT,
  dBusAhb_HRESP,
  iBusAhb_HRDATA,
  iBusAhb_HREADY,
  iBusAhb_HRESP,
  CORE_TDO,
  SYS_RST_o,
  dBusAhb_HADDR,
  dBusAhb_HBURST,
  dBusAhb_HPROT,
  dBusAhb_HREADY_IN,
  dBusAhb_HSIZE,
  dBusAhb_HTRANS,
  dBusAhb_HWDATA,
  dBusAhb_HWRITE,
  dBusAhb_SEL,
  iBusAhb_HADDR,
  iBusAhb_HBURST,
  iBusAhb_HPROT,
  iBusAhb_HSIZE,
  iBusAhb_HTRANS,
  iBusAhb_HWDATA,
  iBusAhb_HWRITE
  );

  input CORE_TCK;
  input CORE_TDI;
  input CORE_TMS;
  input [5:0] INTERRUPT_i;
  input POR_RST_i;
  input SYS_CLK;
  input TIM_CLK;
  input [31:0] dBusAhb_HRDATA;
  input dBusAhb_HREADY_OUT;
  input dBusAhb_HRESP;
  input [31:0] iBusAhb_HRDATA;
  input iBusAhb_HREADY;
  input iBusAhb_HRESP;
  output CORE_TDO;
  output SYS_RST_o;
  output [31:0] dBusAhb_HADDR;
  output [2:0] dBusAhb_HBURST;
  output [3:0] dBusAhb_HPROT;
  output dBusAhb_HREADY_IN;
  output [2:0] dBusAhb_HSIZE;
  output [1:0] dBusAhb_HTRANS;
  output [31:0] dBusAhb_HWDATA;
  output dBusAhb_HWRITE;
  output dBusAhb_SEL;
  output [31:0] iBusAhb_HADDR;
  output [2:0] iBusAhb_HBURST;
  output [3:0] iBusAhb_HPROT;
  output [2:0] iBusAhb_HSIZE;
  output [1:0] iBusAhb_HTRANS;
  output [31:0] iBusAhb_HWDATA;
  output iBusAhb_HWRITE;

  parameter CLSIC_BASEADDR = 16'b0001000000000000;
  parameter CORE_TYPE = "MEDIUM";
  parameter INT_NUM = 6;
  parameter TIC_MTIME_SEL = 1'b0;
  wire [31:0] al_7c5dfaf6;
  wire [5:0] al_d264c8ee;
  wire [5:0] al_f92bb470;
  wire [31:0] al_ad9a3ca4;
  wire [29:0] al_65949b4f;
  wire [29:0] al_eb4cb082;
  wire [29:0] al_831101f2;
  wire [0:0] al_384c501e;
  wire [5:0] al_e108f0ff;
  wire [31:0] al_5d92ff7c;
  wire [3:0] al_5d13c933;
  wire [3:0] al_24e92378;
  wire [31:0] al_45e5d9f7;
  wire [31:0] al_3dcca8e;
  wire [31:0] al_4d9a3d8e;
  wire [3:0] al_7b80e496;
  wire [3:0] al_9d1d880c;
  wire [3:0] al_86d3f01a;
  wire [3:0] al_1a8c7c22;
  wire [31:0] al_ccabc055;
  wire [31:0] al_c28c3a52;
  wire [1:0] al_12792818;
  wire [1:0] al_591b5570;
  wire [31:0] al_97943858;
  wire [29:0] al_35d85285;
  wire [1:0] al_41e76523;
  wire [31:0] al_43722bf9;
  wire [31:0] al_d610ac57;
  wire [4:0] al_6a6a2b33;
  wire [31:0] al_4fd032af;
  wire [31:0] al_8c9327d6;
  wire [31:0] al_40185430;
  wire [31:0] al_a16ef20a;
  wire [30:0] al_b24d99c7;
  wire [31:0] al_bde0dc95;
  wire [15:0] al_5fd02584;
  wire [31:0] al_8778492e;
  wire [31:0] al_f65e6902;
  wire [31:0] al_c1211126;
  wire [31:0] al_126b3afd;
  wire [29:0] al_683f5875;
  wire [2:0] al_9b5530fd;
  wire [31:0] al_adeed2de /* synthesis keep=true */ ;
  wire [32:0] al_b86dd14b;
  wire [31:0] al_cf18c1c6;
  wire [2:0] al_202f2c67;
  wire [2:0] al_b537d840;
  wire [2:0] al_2978b178;
  wire [31:0] al_3bdbe1c8;
  wire [2:0] al_6515336d;
  wire [31:0] al_85a2bdb0;
  wire [31:0] al_1f3eaa15;
  wire [31:0] al_81a1940d;
  wire [31:0] al_8c7f68e2;
  wire [31:0] al_fe073fc9;
  wire [31:0] al_8492e16;
  wire [0:0] al_de0f70d9;
  wire [0:0] al_c50e70c2;
  wire [0:0] al_bb2524be;
  wire [0:0] al_c52295d9;
  wire [0:0] al_4ab1b7b3;
  wire [0:0] al_40dcfa8c;
  wire [0:0] al_361dafb5;
  wire [21:0] al_c6966291;
  wire [0:0] al_192b30b5;
  wire [11:0] al_4a753b95;
  wire [31:0] al_6e268dd3;
  wire [30:0] al_40a6f08c;
  wire [31:0] al_8221e5ce;
  wire [31:0] al_8aeaa5c1;
  wire [31:0] al_192eeeac;
  wire [31:0] al_6fd79ca;
  wire [32:0] al_9e82589f;
  wire [32:0] al_ee1342f7;
  wire [31:0] al_18077581;
  wire [31:0] al_3ca44efd;
  wire [31:0] al_f2330f79;
  wire [31:0] al_94f1da4c;
  wire [32:0] al_32172a12;
  wire [31:0] al_f3b8f942;
  wire [35:0] al_8f26ae38;
  wire [36:1] al_8b049eb2;
  wire [36:1] al_468d3b3e;
  wire [37:0] al_8dd2d746;
  wire [2:0] al_c3eb1e82;
  wire [31:0] al_2cbb16b4;
  wire [31:0] al_8c4e5d9c;
  wire [31:0] al_704d20e3;
  wire [31:0] al_bbc99cd7;
  wire [31:0] al_52ea52d7;
  wire [1:0] al_bb6625de;
  wire [1:0] al_1edb758f;
  wire [1:0] al_580ff8b7;
  wire [1:0] al_b5f1afb5;
  wire [31:0] al_e03b3126;
  wire [31:0] al_9bf95cff;
  wire [31:0] al_8074bdb;
  wire [31:0] al_2f7928e2;
  wire [1:0] al_27c2eb8;
  wire [1:0] al_555b0990;
  wire [1:0] al_a1e88c0c;
  wire [31:0] al_6f2fa5dc;
  wire [31:0] al_d57349d9;
  wire [31:0] al_35295e0a;
  wire [16:0] al_da34572b;
  wire [16:0] al_65e3dd93;
  wire [31:0] al_3e08733b /* synthesis keep=true */ ;
  wire [31:0] al_b541ca02 /* synthesis keep=true */ ;
  wire [31:0] al_46ea2d9f;
  wire [1:0] al_53188262;
  wire [31:0] al_a0e6869c;
  wire [1:0] al_50f87e49;
  wire [33:0] al_3d2fbc2e;
  wire [33:0] al_9edb1d1e;
  wire [31:0] al_ccb50b3a;
  wire [31:0] al_2e7cde15;
  wire [31:0] al_bfc96350;
  wire [1:0] al_727d2e98;
  wire [31:0] al_d1fb6e0a;
  wire [3:0] al_53f57cc3;
  wire [31:0] al_a550c05f;
  wire [33:0] al_d48366e1;
  wire [33:0] al_8eb7c3ef;
  wire [0:0] al_871b264a;
  wire [0:0] al_c2ae0151;
  wire [3:0] al_549b2fd9;
  wire [3:0] al_a3de3eda;
  wire [3:0] al_a6bbd516;
  wire  al_fa675d9c;
  wire [31:0] al_156dfeae;
  wire [4:0] al_cac83419;
  wire [31:0] al_63edc714;
  wire [64:0] al_7b59c46e;
  wire [5:0] al_1d392f4f;
  wire [5:0] al_2d4f70b0;
  wire [31:0] al_ec26021c;
  wire [31:0] al_830b3656;
  wire [32:0] al_a5f7e6c;
  wire [32:0] al_b70cb9be;
  wire [32:0] al_d0c02c51;
  wire [32:0] al_afda7fe3;
  wire [32:0] al_439698e9;
  wire [31:0] al_f12834e3;
  wire [31:0] al_f337bb3c;
  wire [31:0] al_4e7a070d;
  wire [1:0] al_212ac3ba;
  wire [31:0] al_36a894af;
  wire [1:0] al_70c1ae82;
  wire [31:0] al_24ce3017;
  wire [33:0] al_1d8f7667;
  wire [31:0] al_d7ecfd18;
  wire [51:0] al_71c7f8f0;
  wire [31:0] al_e45b51d9;
  wire [31:0] al_8900fb4e;
  wire [44:0] al_de2ed994;
  wire [3:0] al_f1e7f5b0;
  wire [53:0] al_193295bb;
  wire [3:0] al_74afebb7;
  wire [44:0] al_9aa9386d;
  wire [53:0] al_25ac6d54;
  wire [44:0] al_1ee074c7;
  wire [53:0] al_63395efb;
  wire [3:0] al_d4e9c8e0;
  wire [44:0] al_8ffa2af5;
  wire [53:0] al_186e4c3b;
  wire [3:0] al_574e0a5c;
  wire [44:0] al_3d954d6;
  wire [53:0] al_4dc1fe7;
  wire [3:0] al_e1be9e86;
  wire  al_b380555;
  wire [31:0] al_7aa9f4ee;
  wire [31:0] al_f4b0c1c2;
  wire [2:0] al_5c72a609;
  wire [2:0] al_74dc1091;
  wire [2:0] al_a7b01c14;
  wire [2:0] al_fe97bdd9;
  wire [66:0] al_25fbce42;
  wire [7:0] al_8a4a038;
  wire [31:0] al_daece8d7;
  wire al_afa99249;
  wire al_63842eca;
  wire al_aabf3e05;
  wire al_ce484726;
  wire al_6a01eacd;
  wire al_9ab3fa7e;
  wire al_45a5e4cd;
  wire al_5fde6364;
  wire al_98083b2a;
  wire al_b935f70;
  wire al_72cf4613;
  wire al_65e27d78;
  wire al_33785de1;
  wire al_a50da65e;
  wire al_caba2fac;
  wire al_82b381ff;
  wire al_33365b48;
  wire al_c2fc5aeb;
  wire al_6ab36ff1;
  wire al_dd2f78da;
  wire al_8179cfdf;
  wire al_45cc89d;
  wire al_7568a715;
  wire al_4609cf3c;
  wire al_e181a464;
  wire al_b1593081;
  wire al_50a1040b;
  wire al_3e563e21;
  wire al_899000eb;
  wire al_1c92cde;
  wire al_e846ab0b;
  wire al_78f1e056;
  wire al_7704555;
  wire al_6a3d23ee;
  wire al_cffac9df;
  wire al_932f8140;
  wire al_fa1d7661;
  wire al_6f8c3f2d;
  wire al_917164b4;
  wire al_5ce11e05;
  wire al_99e052bc;
  wire al_e84a0f1e;
  wire al_8f7c15b2;
  wire al_133c9e7c;
  wire al_c71e5d62;
  wire al_a2c0d252;
  wire al_9bc5b10b;
  wire al_1df2c985;
  wire al_a99e75eb;
  wire al_7ee9f8d;
  wire al_bd909ea1;
  wire al_80b19a9e;
  wire al_be111ebc;
  wire al_69da6feb;
  wire al_942fb5b3;
  wire al_31800d3e;
  wire al_68c8085f;
  wire al_7a9d9124;
  wire al_e85a2cb7;
  wire al_ccef9e4c;
  wire al_2e06c46d;
  wire al_dc5ae5dc;
  wire al_2fcd16aa;
  wire al_82aaac97;
  wire al_dca31e55;
  wire al_1cf6c96;
  wire al_a4a54bdd;
  wire al_4aafd23e;
  wire al_36b19484;
  wire al_3e310318;
  wire al_a7747a86;
  wire al_ece70a8c;
  wire al_c0f2d5f7;
  wire al_921bc4ca;
  wire al_92eee380;
  wire al_9c367b3e;
  wire al_747f0d5b;
  wire al_4c590039;
  wire al_70d8b4ee;
  wire al_9eda716;
  wire al_29632809;
  wire al_e9c55e9a;
  wire al_4989df73;
  wire al_c3006fde;
  wire al_2c4c1ef7;
  wire al_f325673f;
  wire al_3d3aa49b;
  wire al_8e7f80da;
  wire al_5bcb7210;
  wire al_e2d7fc47;
  wire al_a0b8db17;
  wire al_6f14f6e5;
  wire al_4fdb397d;
  wire al_2672f5b2;
  wire al_82ca9a92;
  wire al_879c97c5;
  wire al_837e8da8;
  wire al_9c95e435;
  wire al_542d1ba4;
  wire al_f4e939bc;
  wire al_26903ef3;
  wire al_82a77528;
  wire al_5b477973;
  wire al_12fa803d;
  wire al_6426fa0c;
  wire al_8b1fccb;
  wire al_4e576557;
  wire al_6c384295;
  wire al_63a3bec2;
  wire al_4a1a4a4;
  wire al_7f54ca49;
  wire al_16541a17;
  wire al_2bfbeb6;
  wire al_1f8435f6;
  wire al_24d740cb;
  wire al_f2f80319;
  wire al_80daf3e;
  wire al_f50ab810;
  wire al_3d0077da;
  wire al_73502252;
  wire al_df3a7245;
  wire al_829d1309;
  wire al_966d08ce;
  wire al_d8039a59;
  wire al_d81efc87;
  wire al_afa2ef7a;
  wire al_5a473143;
  wire al_9a380597;
  wire al_2fd5db25;
  wire al_83abb1fc;
  wire al_bb6e1564;
  wire al_76d86d60;
  wire al_abafb840;
  wire al_665b60c1;
  wire al_9367b2dc;
  wire al_e6c5dfa;
  wire al_5188e109;
  wire al_75b52645;
  wire al_20769005;
  wire al_4d3a4f57;
  wire al_ead254a9;
  wire al_bdce010d;
  wire al_8cc085cf;
  wire al_83e5bc67;
  wire al_cc21f874;
  wire al_304a2593;
  wire al_de514d5;
  wire al_3178c29a;
  wire al_bf8b5005;
  wire al_322e0ef8;
  wire al_9cc77063;
  wire al_5c37ca50;
  wire al_7e8c6cca;
  wire al_1b896d0b;
  wire al_a8c77bd0;
  wire al_3d1aa152;
  wire al_8bea08a7;
  wire al_e9d567fe;
  wire al_bec39e4d;
  wire al_e379ebb5;
  wire al_f6cd735f;
  wire al_c91705db;
  wire al_ea2eaeb1;
  wire al_9d63e9cd;
  wire al_68b106c6;
  wire al_6ec8afa5;
  wire al_2f23ede9;
  wire al_689ac380;
  wire al_17050ddb;
  wire al_6faa66d6;
  wire al_c6d62120;
  wire al_2e313516;
  wire al_2f2822d8;
  wire al_99aa8cdf;
  wire al_2a7e21ae;
  wire al_26f3954d;
  wire al_e4d5d147;
  wire al_c0f96426;
  wire al_8b7c83a7;
  wire al_95a8aeaf;
  wire al_4be831c2;
  wire al_277cf2f2;
  wire al_8ac7c093;
  wire al_c76629d2;
  wire al_a3a8b68d;
  wire al_11418f51;
  wire al_f170970d;
  wire al_c85db05d;
  wire al_a5849610;
  wire al_12227f77;
  wire al_c572d1c7;
  wire al_6a0e908c;
  wire al_c795a432;
  wire al_c197c567;
  wire al_2c3e73df;
  wire al_291d5f8b;
  wire al_cdfe2d97;
  wire al_71fb98b4;
  wire al_5e60a110;
  wire al_4f6deaed;
  wire al_3e5baa1a;
  wire al_134ffa88;
  wire al_33a34bec;
  wire al_6f08d701;
  wire al_dc5d601;
  wire al_39d0a986;
  wire al_fccc3291;
  wire al_37a2cec8;
  wire al_c46301d;
  wire al_f76e538f;
  wire al_b279136c;
  wire al_e0005a94;
  wire al_523a156f;
  wire al_6e8514b8;
  wire al_6a6f79fc;
  wire al_7daf5294;
  wire al_cc4ef047;
  wire al_e9183b70;
  wire al_7709e0b8;
  wire al_5907d462;
  wire al_e83c9381;
  wire al_b4c2dbf;
  wire al_cd728703;
  wire al_6dc2ee9d;
  wire al_36d94dee;
  wire al_e493cfe2;
  wire al_a122473;
  wire al_571b50e9;
  wire al_91e1bb2e;
  wire al_89941f61;
  wire al_57355198;
  wire al_c768664c;
  wire al_7e44038b;
  wire al_c6e3e50;
  wire al_58a3b7ac;
  wire al_fe608411;
  wire al_a8c327eb;
  wire al_c02355f;
  wire al_50f055e6;
  wire al_7971debc;
  wire al_8628bcb0;
  wire al_5d524bff;
  wire al_ed4da032;
  wire al_931aa04b;
  wire al_571c1ade;
  wire al_7d44614a;
  wire al_fc020630;
  wire al_381491bf;
  wire al_862095a3;
  wire al_4348da93;
  wire al_3c0b578d;
  wire al_8c1979b0;
  wire al_6a1d2e79;
  wire al_1520e815;
  wire al_7bc70fec;
  wire al_5b63e1bd;
  wire al_c30b4452;
  wire al_1da1b47c;
  wire al_f380f225;
  wire al_c45763da;
  wire al_91dd025b;
  wire al_1e473c0d;
  wire al_429b8bb;
  wire al_a0d06894;
  wire al_ab3758ac;
  wire al_399d7ca4;
  wire al_e87887db;
  wire al_252ad8ef;
  wire al_ed00e897;
  wire al_5ab03ac;
  wire al_6afd474a;
  wire al_ae709366;
  wire al_1a6b06a2;
  wire al_630fb1c3;
  wire al_ac5e9239;
  wire al_f58e845f;
  wire al_388498bb;
  wire al_9ef79df4;
  wire al_818b914;
  wire al_b113fb3b;
  wire al_614db1c3;
  wire al_8dd6f665;
  wire al_2340ada;
  wire al_6233890d;
  wire al_d0d487f0;
  wire al_f5ef5e84;
  wire al_dea86dcd;
  wire al_429d51be;
  wire al_c5f16127;
  wire al_9b8294d5;
  wire al_382bcd96;
  wire al_59258acc;
  wire al_5a3cd9;
  wire al_e3fa7139;
  wire al_a4b5d1d0;
  wire al_774d209c;
  wire al_eecd0df4;
  wire al_491245fc;
  wire al_151b9283;
  wire al_aac49860;
  wire al_826899ea;
  wire al_3401493;
  wire al_e381eae8;
  wire al_29590532;
  wire al_a5dcf577;
  wire al_f20e1999;
  wire al_9f91dd62;
  wire al_4945d0da;
  wire al_7cba307c;
  wire al_50fdf48e;
  wire al_bc2094a;
  wire al_be7d7ec3;
  wire al_7c4abb1c;
  wire al_35216c23;
  wire al_34eb7e40;
  wire al_8bbc936e;
  wire al_33f7e9f;
  wire al_82cf60b4;
  wire al_87a252af;
  wire al_e2de4855;
  wire al_6e34d4cd;
  wire al_1af3cc59;
  wire al_2161900e;
  wire al_eba13280;
  wire al_837ccd29;
  wire al_9711882c;
  wire al_2d65cded;
  wire al_de77c599;
  wire al_e2f41361;
  wire al_af2b71d8;
  wire al_96191e5;
  wire al_b81cc851;
  wire al_1af8f97e;
  wire al_4db67ec5;
  wire al_24887a1a;
  wire al_9a21e871;
  wire al_35d69006;
  wire al_d3f03020;
  wire al_2d292595;
  wire al_5325cd47;
  wire al_bf79dcf1;
  wire al_58ec462a;
  wire al_42d8598b;
  wire al_9bb4d4a4;
  wire al_82229532;
  wire al_ec42a4de;
  wire al_4aed8be6;
  wire al_9cf531f8;
  wire al_a430e4d2;
  wire al_98ab69b8;
  wire al_5f3d7b85;
  wire al_1b14c7a0;
  wire al_fc39fece;
  wire al_d1df0873;
  wire al_b4eb77a8;
  wire al_4ed9ad89;
  wire al_955e8db5;
  wire al_22883704;
  wire al_3f04848f;
  wire al_6c5ae138;
  wire al_89ab45b5;
  wire al_2dc65bff;
  wire al_2c78771b;
  wire al_271667bb;
  wire al_25ff0fe3;
  wire al_d3323cee;
  wire al_6be7ae97;
  wire al_c2ce02d3;
  wire al_fdcd8a4d;
  wire al_92a03ec7;
  wire al_72cf1502;
  wire al_53cc722d;
  wire al_c85e3cfa;
  wire al_695857c1;
  wire al_583b2c0d;
  wire al_73767b69;
  wire al_22240f9f;
  wire al_e9e54e67;
  wire al_dfe2f2a3;
  wire al_dbe911b7;
  wire al_a7fbaeb;
  wire al_59bca917;
  wire al_c92e4639;
  wire al_a5d442e7;
  wire al_91974942;
  wire al_d135ca94;
  wire al_ab9e30a4;
  wire al_4d279efb;
  wire al_ae1b5d59;
  wire al_f466006e;
  wire al_4d64c75;
  wire al_5a617f02;
  wire al_c63a3306;
  wire al_6b46d3b9;
  wire al_8c8f6789;
  wire al_443b56a1;
  wire al_19286ed8;
  wire al_82a462e4;
  wire al_2f093a42;
  wire al_debb551a;
  wire al_cd5a3103;
  wire al_24003c83;
  wire al_ec08a0e6;
  wire al_c06b4d62;
  wire al_c862b555;
  wire al_c28f9c66;
  wire al_3f573e25;
  wire al_62997e0b;
  wire al_6076534a;
  wire al_5e07bd5e;
  wire al_4efe0c98;
  wire al_c64cf9f6;
  wire al_89bb053a;
  wire al_ecd761fc;
  wire al_a155e0b3;
  wire al_9852e0df;
  wire al_193c583f;
  wire al_f19f190e;
  wire al_ad2a00e5;
  wire al_debfa536;
  wire al_faaecf2;
  wire al_267d2aa;
  wire al_89782fa0;
  wire al_5ca98598;
  wire al_40d63aa3;
  wire al_f814979a;
  wire al_5a93aea7;
  wire al_6758eae2;
  wire al_42b103ed;
  wire al_e2259475;
  wire al_b40171bd;
  wire al_82b168eb;
  wire al_20b06ef3;
  wire al_89a93b84;
  wire al_b6803a27;
  wire al_2eb5050b;
  wire al_7bf844c2;
  wire al_d0702be9;
  wire al_afd990ff;
  wire al_f5f3edb6;
  wire al_9df5b848;
  wire al_5b3ba944;
  wire al_d1fc8906;
  wire al_2fb7633;
  wire al_afe5948f;
  wire al_2d354b;
  wire al_be6e0599;
  wire al_c89d1229;
  wire al_1953385a;
  wire al_70f172be;
  wire al_cc989ac9;
  wire al_8d9bdfff;
  wire al_2cd19c12;
  wire al_a89113a9;
  wire al_e3fa27d;
  wire al_fd8d8e0c;
  wire al_7b4ebd2a;
  wire al_6ab73d4d;
  wire al_c585508d;
  wire al_63bbd3a2;
  wire al_45322fba;
  wire al_263322e4;
  wire al_22da7862;
  wire al_a3f3ee06;
  wire al_3ab03292;
  wire al_428b50b6;
  wire al_5bcd7a0;
  wire al_ca581e6c;
  wire al_cc5bfca5;
  wire al_e79b3dfa;
  wire al_6ae2a07d;
  wire al_4d016a39;
  wire al_14b732b9;
  wire al_cacb44c4;
  wire al_19c0990d;
  wire al_cae21d2e;
  wire al_d78f6bd4;
  wire al_a69cec28;
  wire al_9b707062;
  wire al_3a7c5a5;
  wire al_2ede456b;
  wire al_bf6a3977;
  wire al_30f08f9c;
  wire al_3656d228;
  wire al_cd498e9f;
  wire al_f430a5aa;
  wire al_eead7739;
  wire al_5727b773;
  wire al_8488923;
  wire al_59be2ab1;
  wire al_c8ba6c61;
  wire al_b5bf2603;
  wire al_fdf9f0dc;
  wire al_407c8ac1;
  wire al_728c73ac;
  wire al_a35cf148;
  wire al_a6e0ed04;
  wire al_e163f204;
  wire al_8e267e24;
  wire al_5df930ee;
  wire al_1e979a01;
  wire al_80e2c141;
  wire al_512b1421;
  wire al_1891b3c7;
  wire al_60dd36d7;
  wire al_f1bb92e9;
  wire al_3626cb0;
  wire al_3b8c31d7;
  wire al_102b7ad2;
  wire al_6ec45564;
  wire al_e611ec68;
  wire al_53b3dbc6;
  wire al_1f5093b5;
  wire al_ffc4fe26;
  wire al_658bb789;
  wire al_a831c176;
  wire al_c7df4b4d;
  wire al_3b0f4da7;
  wire al_d76255c5;
  wire al_7d27d680;
  wire al_f61ec828;
  wire al_7e6320f4;
  wire al_e6455839;
  wire al_d00a6f56;
  wire al_3ebb68c3;
  wire al_98804c07;
  wire al_6d92b3c6;
  wire al_bdb28b76;
  wire al_73fb1ee5;
  wire al_33a2911e;
  wire al_8a841cb4;
  wire al_c861c8f0;
  wire al_76a52f3d;
  wire al_bf952132;
  wire al_2370214;
  wire al_f4b5275b;
  wire al_e5ffe4ff;
  wire al_36d679eb;
  wire al_ce0d355f;
  wire al_bd56460d;
  wire al_c0406dbc;
  wire al_14651309;
  wire al_730b0315;
  wire al_dc741944;
  wire al_86608ce5;
  wire al_1e27127a;
  wire al_8675b08;
  wire al_f465aa2;
  wire al_79fcc7dd;
  wire al_44ee9376;
  wire al_b6d6e907;
  wire al_f8b84ed9;
  wire al_278217fa;
  wire al_d66e22dd;
  wire al_9ce6f9ae;
  wire al_1b5c5256;
  wire al_bc831201;
  wire al_36303862;
  wire al_569f263c;
  wire al_b1924903;
  wire al_41adb443;
  wire al_b5b0f369;
  wire al_5c3a44f0;
  wire al_3cd3f418;
  wire al_c78a6044;
  wire al_7b2239bb;
  wire al_f2fcadd6;
  wire al_50c53403;
  wire al_289dceb2;
  wire al_dc412458;
  wire al_f0561e92;
  wire al_319b4c4c;
  wire al_10df355f;
  wire al_ed766401;
  wire al_23658752;
  wire al_e9a9157c;
  wire al_7b880725;
  wire al_7750a3cd;
  wire al_70fea121;
  wire al_385f14;
  wire al_bb4f8966;
  wire al_6d174013;
  wire al_14816c03;
  wire al_ce80e68f;
  wire al_dfe3b0a5;
  wire al_cb828215;
  wire al_80b925b7;
  wire al_65a874f0;
  wire al_8a79ceb4;
  wire al_5c0f2717;
  wire al_daaf28b4;
  wire al_bf987e25;
  wire al_b44f8827;
  wire al_f49386;
  wire al_f6c8a5f0;
  wire al_94f9539;
  wire al_5914a559;
  wire al_85bef49;
  wire al_354f5999;
  wire al_92fd4928;
  wire al_29a1a38f;
  wire al_26af78f7;
  wire al_37698acd;
  wire al_bb5767ca;
  wire al_75b09ba0;
  wire al_7095ffb4;
  wire al_e0306332;
  wire al_a34c4405;
  wire al_a0c987d5;
  wire al_bdfc704c;
  wire al_f4418953;
  wire al_193dedee;
  wire al_c0855656;
  wire al_fdd40d67;
  wire al_63c14fc;
  wire al_48dfd35c;
  wire al_1de941c8;
  wire al_5f34afe1;
  wire al_10ccc4a2;
  wire al_7fea1a88;
  wire al_90ed329;
  wire al_6d5a6293;
  wire al_aa88d0b2;
  wire al_6ecad7e7;
  wire al_42d0475;
  wire al_927566f;
  wire al_18e9bd9b;
  wire al_e2f2e915;
  wire al_d0a81721;
  wire al_f529ac86;
  wire al_13bd3caf;
  wire al_52ea8e26;
  wire al_f0a4b18b;
  wire al_1e389db1;
  wire al_123d8e5f;
  wire al_a241616a;
  wire al_8e70d65a;
  wire al_45ceabc3;
  wire al_19e34f5d;
  wire al_9a97f855;
  wire al_edcbe33d;
  wire al_91a72f10;
  wire al_a59daeb4;
  wire al_781bb51f;
  wire al_d4ff0ad3;
  wire al_ffb1962;
  wire al_443f5c3a;
  wire al_d2147867;
  wire al_1e7955bd;
  wire al_9bb19ed8;
  wire al_ac5b8836;
  wire al_ee66e790;
  wire al_1c02d8ab;
  wire al_8db3355a;
  wire al_dd37dc5d;
  wire al_cae3c642;
  wire al_e87ca79;
  wire al_74973e72;
  wire al_a0670bff;
  wire al_447f0158;
  wire al_b62de081;
  wire al_d33dd538;
  wire al_ab46d2b9;
  wire al_825438f5;
  wire al_f76f8d54;
  wire al_6e8dae0d;
  wire al_31822056;
  wire al_c6cd8be8;
  wire al_c048f5a0;
  wire al_c5cc2f9b;
  wire al_8cb8f5f5;
  wire al_13708b94;
  wire al_c4d4b7f5;
  wire al_fb26226a;
  wire al_667db93d;
  wire al_4ed450cb;
  wire al_4a696460;
  wire al_2418b5af;
  wire al_4e819ed5;
  wire al_640ea1c6;
  wire al_8773b31;
  wire al_3be09bce;
  wire al_e9dadc09;
  wire al_3db1ed2d;
  wire al_81e43d4;
  wire al_24cba21e;
  wire al_6cfd8dcf;
  wire al_a2aa312d;
  wire al_5beecaa3;
  wire al_3b6c54b6;
  wire al_50439dee;
  wire al_72de3c0a;
  wire al_b0555243;
  wire al_210b38e6;
  wire al_bbee20b8;
  wire al_c1d3ffb3;
  wire al_3e1875be;
  wire al_27878642;
  wire al_ac867fa2;
  wire al_8b9b5b1d;
  wire al_80a6299b;
  wire al_6305766;
  wire al_e51dc3c;
  wire al_5fe5e97d;
  wire al_35379d79;
  wire al_5a3ca2c7;
  wire al_e791df33;
  wire al_168ce6c3;
  wire al_1e8c20b0;
  wire al_5a6794e3;
  wire al_d3114685;
  wire al_4ea1bb54;
  wire al_d5e048cf;
  wire al_1eaad5d4;
  wire al_c63ed4c6;
  wire al_cd3394ba;
  wire al_b2f6a2a2;
  wire al_b63bb946;
  wire al_abfe390c;
  wire al_da123ab6;
  wire al_f92423e;
  wire al_b9001309;
  wire al_d56de4dc;
  wire al_3e7bf97e;
  wire al_e99a5572;
  wire al_47e27082;
  wire al_ea06ea2d;
  wire al_8b49a361;
  wire al_dccb8299;
  wire al_bd675004;
  wire al_22e7124d;
  wire al_1c537db1;
  wire al_bbb6292e;
  wire al_4c1d95c5;
  wire al_39ff3661;
  wire al_a60ca806;
  wire al_370b9296;
  wire al_3cd3cca9;
  wire al_126b9a65;
  wire al_f57c7577;
  wire al_dffeb202;
  wire al_343c5862;
  wire al_a683a564;
  wire al_57675c9b;
  wire al_997b23f2;
  wire al_f1e867e0;
  wire al_69efc6c6;
  wire al_a8d5d0d5;
  wire al_4df86c43;
  wire al_43099296;
  wire al_c51bf9b;
  wire al_136ceed1;
  wire al_ffe7e6d4;
  wire al_b931d891;
  wire al_1bae5100;
  wire al_8bc7d472;
  wire al_55994c98;
  wire al_2137298d;
  wire al_b0c44f4;
  wire al_da3cc173;
  wire al_c017beac;
  wire al_96f2b26a;
  wire al_d50e9dc4;
  wire al_4c6b15c2;
  wire al_57bbe3ad;
  wire al_f7e849b8;
  wire al_2978bc8a;
  wire al_c8e314e6;
  wire al_f2b407ac;
  wire al_c6dd3893;
  wire al_b4d3ef2b;
  wire al_70eedb8b;
  wire al_d7081cd4;
  wire al_792f120f;
  wire al_77120298;
  wire al_a32b870b;
  wire al_c96d1fd5;
  wire al_479534eb;
  wire al_56afc96e;
  wire al_28a777ae;
  wire al_94dd833a;
  wire al_ba6916cf;
  wire al_357abca7;
  wire al_d2ba0b0;
  wire al_4712f186;
  wire al_8fddd1ab;
  wire al_df5cc0b8;
  wire al_5b3d235a;
  wire al_9a488676;
  wire al_9ae3000c;
  wire al_5c28a20d;
  wire al_8f175a04;
  wire al_349edb3b;
  wire al_c6c291a5;
  wire al_865e8f41;
  wire al_2ac34e44;
  wire al_dfd548fb;
  wire al_90ba8dd5;
  wire al_cee3e376;
  wire al_fb22b66;
  wire al_83a071a4;
  wire al_55ed4df1;
  wire al_f03f7670;
  wire al_dfdc4f07;
  wire al_6df79c7b;
  wire al_7c75aadd;
  wire al_f7b11965;
  wire al_74e1f810;
  wire al_5c743358;
  wire al_87b30ed5;
  wire al_e22f5efa;
  wire al_286b6a5c;
  wire al_d344e0e5;
  wire al_2d35601b;
  wire al_6e7063d6;
  wire al_8647937a;
  wire al_c524b83f;
  wire al_55bbd6fb;
  wire al_7c8ae043;
  wire al_7244a2ec;
  wire al_52be31ea;
  wire al_1dcba582;
  wire al_8906de47;
  wire al_9df643fa;
  wire al_568af2d5;
  wire al_97cb05f;
  wire al_47eda15e;
  wire al_c6ff495c;
  wire al_2f34d7b4;
  wire al_e3502e80;
  wire al_4002af45;
  wire al_77bf7190;
  wire al_843f038d;
  wire al_1f0371f8;
  wire al_31f2e639;
  wire al_ba3f2ea7;
  wire al_7a7cc81;
  wire al_bdf9a7dd;
  wire al_653f9409;
  wire al_3629238d;
  wire al_12584de1;
  wire al_65dc271;
  wire al_f5b7debb;
  wire al_a8af8112;
  wire al_42488c02;
  wire al_af575898;
  wire al_bd10bda8;
  wire al_c7467d2d;
  wire al_e240543c;
  wire al_88a18e08;
  wire al_1754eacf;
  wire al_a72e375d;
  wire al_2df3af97;
  wire al_3f6865d3;
  wire al_3577d7b9;
  wire al_dec34edc;
  wire al_79632d6f;
  wire al_12790a23;
  wire al_c115942c;
  wire al_d68a240f;
  wire al_3ce9d83;
  wire al_19463fbe;
  wire al_ef0a8112;
  wire al_14c6d47a;
  wire al_d63f10c0;
  wire al_9e9618ab;
  wire al_c74661;
  wire al_387eb97;
  wire al_d7a80970;
  wire al_d84a4a58;
  wire al_88242571;
  wire al_ff37bd99;
  wire al_b0110a42;
  wire al_75ee8673;
  wire al_33012db3;
  wire al_b4ed90bc;
  wire al_90d6c009;
  wire al_ec9911d2;
  wire al_ce46ef05;
  wire al_78e2749c;
  wire al_e1adfd34;
  wire al_ac6ff6aa;
  wire al_31e9afe8;
  wire al_575fad37;
  wire al_2a0680fd;
  wire al_c964851;
  wire al_4e9ff654;
  wire al_ea114973;
  wire al_2dba6136;
  wire al_4cc73535;
  wire al_4381d4c9;
  wire al_3c39e4b0;
  wire al_d9533dba;
  wire al_a7a12e87;
  wire al_7daf0c48;
  wire al_fb6b4008;
  wire al_d41aa0e7;
  wire al_a4f54b87;
  wire al_71df23fe;
  wire al_d9a23597;
  wire al_76cdacda;
  wire al_74831af1;
  wire al_97966a28;
  wire al_ae1d4fee;
  wire al_5281bd0f;
  wire al_784638ef;
  wire al_8bfeeae9;
  wire al_f6c0774b;
  wire al_3833a138;
  wire al_fc3546f;
  wire al_c14f8945;
  wire al_3a175d67;
  wire al_6c7e2f3;
  wire al_897eb9f3;
  wire al_efb93bad;
  wire al_de36fb50;
  wire al_4f8cbab6;
  wire al_3c3c44e5;
  wire al_2edab7d3;
  wire al_786d2b97;
  wire al_723a595b;
  wire al_42c07e1a;
  wire al_d6c2acee;
  wire al_dd28d822;
  wire al_be8dbeba;
  wire al_460aa351;
  wire al_18e8ea79;
  wire al_4183cccb;
  wire al_f405df5e;
  wire al_cb204385;
  wire al_fb048e7c;
  wire al_e9d7a836;
  wire al_d1b00369;
  wire al_3789ddb5;
  wire al_30a65d08;
  wire al_9617ef5a;
  wire al_cf16e2e3;
  wire al_8953e749;
  wire al_6c0635b4;
  wire al_1fb1fe24;
  wire al_5a1a38b6;
  wire al_2b49ac1e;
  wire al_9dba4e2f;
  wire al_68b1ca17;
  wire al_286e2d87;
  wire al_7b1d42ce;
  wire al_4bbe4f7c;
  wire al_edead58e;
  wire al_5eff1a16;
  wire al_a860806e;
  wire al_db9a596c;
  wire al_2beb9d89;
  wire al_aae16022;
  wire al_21fa7d09;
  wire al_bfcbc23b;
  wire al_8e2aeac5;
  wire al_cb20b6b1;
  wire al_362ab5dc;
  wire al_b509771d;
  wire al_3813142e;
  wire al_73cede3c;
  wire al_4605c5c6;
  wire al_2bed4baa;
  wire al_deac45a7;
  wire al_819b6344;
  wire al_1ae2d65b;
  wire al_ab419e9c;
  wire al_4db2159c;
  wire al_b0f1a2c;
  wire al_97c3f56c;
  wire al_a3cc9c36;
  wire al_359eb4b6;
  wire al_fa3c0cbe;
  wire al_13e3d996;
  wire al_b67365e0;
  wire al_2444302e;
  wire al_8492fa3d;
  wire al_c82d2f1e;
  wire al_af9af7c7;
  wire al_94d4afd7;
  wire al_cdec8c3f;
  wire al_7d5e05f7;
  wire al_6b6f1ca9;
  wire al_722a720c;
  wire al_eb3feb88;
  wire al_35e93aaa;
  wire al_aca053a7;
  wire al_45d4540c;
  wire al_d71e234e;
  wire al_ad86ef7d;
  wire al_aa329d99;
  wire al_9d940ee8;
  wire al_e4ddc7f7;
  wire al_a9bc0459;
  wire al_893ad164;
  wire al_cae74074;
  wire al_1a1782f2;
  wire al_b184fe5a;
  wire al_cae48ea4;
  wire al_82238017;
  wire al_43aa4702;
  wire al_162afaa8;
  wire al_59035248;
  wire al_177c2401;
  wire al_d2548651;
  wire al_d5e15803;
  wire al_fbf0401d;
  wire al_e8e20039;
  wire al_692e1afb;
  wire al_5bc78df0;
  wire al_541e0d8b;
  wire al_b950f9ad;
  wire al_63f22050;
  wire al_7a187fb8;
  wire al_3386891f;
  wire al_5278baaa;
  wire al_2295e150;
  wire al_bef23915;
  wire al_90adbe55;
  wire al_ed7763f6;
  wire al_1ab00333;
  wire al_3829588f;
  wire al_12251cca;
  wire al_618e5cf5;
  wire al_a7e3ba76;
  wire al_2e8a294f;
  wire al_90b4cab0;
  wire al_f41fca3f;
  wire al_89494e6b;
  wire al_781ea417;
  wire al_21c33d70;
  wire al_ea118cf6;
  wire al_71c814f5;
  wire al_a478b55f;
  wire al_e7747da7;
  wire al_e3773112;
  wire al_de44ed56;
  wire al_18153c5c;
  wire al_89d8e10c;
  wire al_95046a85;
  wire al_16eb3ffd;
  wire al_d358a549;
  wire al_88c7c32a;
  wire al_74b0792c;
  wire al_dea79dda;
  wire al_36f32db5;
  wire al_7989383a;
  wire al_f176a1bb;
  wire al_bee19057;
  wire al_e3e05361;
  wire al_cbe76bf6;
  wire al_1dab850a;
  wire al_3e17171c;
  wire al_9328cdb4;
  wire al_25614342;
  wire al_477e72e5;
  wire al_d2b99696;
  wire al_d6db317;
  wire al_f7851a1a;
  wire al_12004dbe;
  wire al_7fc6feef;
  wire al_406777f2;
  wire al_79961e57;
  wire al_53750577;
  wire al_568ed982;
  wire al_1a113696;
  wire al_51a7aab3;
  wire al_433e30e8;
  wire al_81feda1d;
  wire al_b669e5e6;
  wire al_a8b9ff36;
  wire al_e8448fdd;
  wire al_71cdacfd;
  wire al_467f9b5e;
  wire al_f48cb7f2;
  wire al_d83ea51;
  wire al_93600cc2;
  wire al_63e36edf;
  wire al_495a58bd;
  wire al_26f7099d;
  wire al_972ccb4f;
  wire al_bd6aed53;
  wire al_ba428019;
  wire al_18cae8b9;
  wire al_92bdd050;
  wire al_cb40733a;
  wire al_428c2665;
  wire al_77af043a;
  wire al_c99791ac;
  wire al_18a866ae;
  wire al_9cb94e30;
  wire al_1e7370cf;
  wire al_1712bb7c;
  wire al_3043d922;
  wire al_69790d6e;
  wire al_b1c0d1f7;
  wire al_58533fed;
  wire al_fa53107d;
  wire al_7a87cf81;
  wire al_3ca77acd;
  wire al_19663434;
  wire al_8e3e7ef7;
  wire al_1df72327;
  wire al_f07170fc;
  wire al_5632987e;
  wire al_c5c038e7;
  wire al_e56ae954;
  wire al_83a5fe89;
  wire al_ad72d731;
  wire al_e6ba0c27;
  wire al_41cca93a;
  wire al_19790099;
  wire al_ab63694b;
  wire al_35ca4317;
  wire al_32a84555;
  wire al_9b78efe2;
  wire al_4507eb5c;
  wire al_627e0d7d;
  wire al_f036124a;
  wire al_6291136b;
  wire al_a27f756f;
  wire al_c4074784;
  wire al_7d2c853e;
  wire al_5fe8f9ad;
  wire al_b469f7cc;
  wire al_9a3c3a5;
  wire al_d508bbc9;
  wire al_d79e66b7;
  wire al_6499e5fd;
  wire al_5e3d90d7;
  wire al_66ffb9;
  wire al_119831c0;
  wire al_5e275e81;
  wire al_b567677b;
  wire al_c871f2ad;
  wire al_4d82afcf;
  wire al_ee8b2558;
  wire al_da7f07ab;
  wire al_aa37cfdb;
  wire al_172eec6a;
  wire al_8869249d;
  wire al_3697c94f;
  wire al_8de27684;
  wire al_a1a600b6;
  wire al_ac1a4f11;
  wire al_74d8fce0;
  wire al_7b361041;
  wire al_3d3ab166;
  wire al_1d8052bb;
  wire al_4d792cee;
  wire al_c1679159;
  wire al_1b41bac1;
  wire al_7242df1f;
  wire al_83268b9b;
  wire al_16745a5f;
  wire al_a63110e1;
  wire al_f5b6a552;
  wire al_75e66ec7;
  wire al_2a43721c;
  wire al_d119a42b;
  wire al_afb86315;
  wire al_67635cb3;
  wire al_8c0460e8;
  wire al_76e89bee;
  wire al_6893b11d;
  wire al_30c029d2;
  wire al_2482626f;
  wire al_6f63d541;
  wire al_8805aafa;
  wire al_52c6af0a;
  wire al_8f2c85dc;
  wire al_b799bc04;
  wire al_50debbc6;
  wire al_69807e37;
  wire al_ddfd7daa;
  wire al_f66ced67;
  wire al_b3a31b1c;
  wire al_48d2ef94;
  wire al_7408b2ea;
  wire al_6897cc6d;
  wire al_766b3b75;
  wire al_da9c21fb;
  wire al_d72f4570;
  wire al_bccf82af;
  wire al_f56de171;
  wire al_e72a5b80;
  wire al_d485b6de;
  wire al_2d6e7982;
  wire al_a2250ee;
  wire al_9c16c2f5;
  wire al_61085a1a;
  wire al_f0ecd262;
  wire al_519869c;
  wire al_536fd7fd;
  wire al_fa66b6a3;
  wire al_bd9d7d67;
  wire al_a25a6119;
  wire al_8c22c3eb;
  wire al_cc14dad7;
  wire al_4bfb7d3a;
  wire al_bcf22cd5;
  wire al_96c3cafb;
  wire al_2cce4860;
  wire al_420d5318;
  wire al_383f9835;
  wire al_1405651f;
  wire al_a40c439;
  wire al_de666865;
  wire al_4cc97ac1;
  wire al_1d7074bf;
  wire al_7a486383;
  wire al_3d334d88;
  wire al_a2deaa78;
  wire al_fa0903ac;
  wire al_f49992c3;
  wire al_94c23c7d;
  wire al_24a3e858;
  wire al_c73c0ba3;
  wire al_b3684022;
  wire al_b8437eb4;
  wire al_eb46e9d2;
  wire al_a8c60ee7;
  wire al_9ba628cf;
  wire al_118827bc;
  wire al_66fb6e33;
  wire al_17dd8854;
  wire al_d5b6b580;
  wire al_b8ccdc1c;
  wire al_84a0e6;
  wire al_c0c7b1b4;
  wire al_acac884e;
  wire al_d020f13b;
  wire al_3d9557e1;
  wire al_628a9731;
  wire al_13f338be;
  wire al_f9c1044d;
  wire al_2c5a98b1;
  wire al_2d4bf1ba;
  wire al_a840afb1;
  wire al_220ba3d7;
  wire al_95cc331e;
  wire al_69c28a29;
  wire al_e92fad27;
  wire al_61365560;
  wire al_5b8651b5;
  wire al_660ff49e;
  wire al_5824822d;
  wire al_951b8fda;
  wire al_6d9a66ce;
  wire al_87fbe8d;
  wire al_8f3d3123;
  wire al_1b1495c6;
  wire al_39f4f94a;
  wire al_9ba605ab;
  wire al_a7eb7455;
  wire al_ac27d20b;
  wire al_271d0926;
  wire al_48e8a022;
  wire al_c21c784f;
  wire al_ac17e182;
  wire al_28aac2f6;
  wire al_bdd9239c;
  wire al_d14a1180;
  wire al_470c29ce;
  wire al_7ba3de08;
  wire al_99df9c8d;
  wire al_7428b0ee;
  wire al_7b0b987;
  wire al_5d89de3c;
  wire al_fb1aae;
  wire al_b8cddd4;
  wire al_8a026941;
  wire al_20e2d49e;
  wire al_5fe9efd2;
  wire al_68a3d338;
  wire al_a4f21dd7;
  wire al_589bdcdb;
  wire al_c83b3308;
  wire al_698ba8c2;
  wire al_ba08f61a;
  wire al_a8151162;
  wire al_b8fe1a1f;
  wire al_d4a46bf1;
  wire al_1a09507b;
  wire al_681bbb63;
  wire al_510fa565;
  wire al_4cb17b0d;
  wire al_566f1754;
  wire al_2434efda;
  wire al_c4aa9af;
  wire al_5978317;
  wire al_170fdda;
  wire al_3f1d46e5;
  wire al_ebace85;
  wire al_6b2d5c80;
  wire al_6715e869;
  wire al_39cb3b56;
  wire al_cbdc72d2;
  wire al_8bf5da64;
  wire al_c5b8f9ea;
  wire al_9a05e7eb;
  wire al_3e46fbe7;
  wire al_9bcd349b;
  wire al_32fedef4;
  wire al_86fb87b9;
  wire al_44595135;
  wire al_36962d69;
  wire al_aded6184;
  wire al_df7b4407;
  wire al_7bc36116;
  wire al_4357844d;
  wire al_eebab250;
  wire al_e2608c20;
  wire al_168e1cf3;
  wire al_2c27d715;
  wire al_6631dfe9;
  wire al_f3435a5b;
  wire al_cdd52893;
  wire al_626d1d9f;
  wire al_ad3403a8;
  wire al_faa08495;
  wire al_4580e6f4;
  wire al_5b3bb87e;
  wire al_5c333c82;
  wire al_8e80a953;
  wire al_43f03d72;
  wire al_13e18942;
  wire al_bdade024;
  wire al_235de557;
  wire al_82a1cc96;
  wire al_c36f1efd;
  wire al_6f3fdf2e;
  wire al_e9897485;
  wire al_163b1f63;
  wire al_9c55c5c3;
  wire al_dc7b4f80;
  wire al_804ebeec;
  wire al_49e80206;
  wire al_d19b9f6b;
  wire al_4bc88254;
  wire al_c281f5b2;
  wire al_be8ea5e1;
  wire al_6782a2e8;
  wire al_4cc0b8dd;
  wire al_58fb1503;
  wire al_7610b7fc;
  wire al_895aceff;
  wire al_a4b1734c;
  wire al_d26be51c;
  wire al_809b319;
  wire al_709aaff2;
  wire al_bb6ca07d;
  wire al_cf7a2555;
  wire al_9176d089;
  wire al_a994b7f;
  wire al_592c9a6;
  wire al_5a744f0f;
  wire al_523cde28;
  wire al_7c88a272;
  wire al_673a4598;
  wire al_cd3d5e6f;
  wire al_cdace779;
  wire al_b2739b77;
  wire al_e3290619;
  wire al_e3edcf1a;
  wire al_587b9831;
  wire al_24641d37;
  wire al_abe3d564;
  wire al_691a2d0a;
  wire al_4f8cc1b7;
  wire al_f36bf4fd;
  wire al_9526c852;
  wire al_a167c8cf;
  wire al_86466d94;
  wire al_76ffd29c;
  wire al_def94157;
  wire al_62da7380;
  wire al_524d11ae;
  wire al_eddc4d82;
  wire al_84c23d54;
  wire al_b968fef9;
  wire al_98842338;
  wire al_bb0cd305;
  wire al_1a1af7e4;
  wire al_501dbbdf;
  wire al_82faef35;
  wire al_41e75372;
  wire al_2af4b91;
  wire al_1ca0e00e;
  wire al_b211b12d;
  wire al_1d840c32;
  wire al_e4d248a4;
  wire al_3f2c3141;
  wire al_8905c135;
  wire al_6f809586;
  wire al_1d3bfd2e;
  wire al_7167debf;
  wire al_5493f072;
  wire al_a2426a1;
  wire al_a62203af;
  wire al_df2df2f9;
  wire al_358f5bea;
  wire al_a559a13b;
  wire al_99763382;
  wire al_1a551855;
  wire al_c0a7a5f;
  wire al_a96ccffb;
  wire al_2b6037c7;
  wire al_acd38e8e;
  wire al_4736f54a;
  wire al_d518b626;
  wire al_5c1a51fa;
  wire al_ab1643c6;
  wire al_bc4322fc;
  wire al_c3666229;
  wire al_d9ff9b46;
  wire al_9061aac4;
  wire al_ac066a39;
  wire al_3d575f81;
  wire al_d72457d3;
  wire al_ee5ae3ff;
  wire al_45c565e6;
  wire al_fbb53e44;
  wire al_a44ada9e;
  wire al_2802ceac;
  wire al_f5a4c6e6;
  wire al_56c9e07a;
  wire al_a4860493;
  wire al_a45b58d1;
  wire al_8bf04ef0;
  wire al_b7e97af1;
  wire al_4c35eef2;
  wire al_59c9e271;
  wire al_31e2d17a;
  wire al_d7a8be80;
  wire al_13a562ab;
  wire al_b5356e8f;
  wire al_6380dbe7;
  wire al_e7b5abb5;
  wire al_c4f8cd6c;
  wire al_53ca6362;
  wire al_6d28932f;
  wire al_eeed7a72;
  wire al_38acf7c0;
  wire al_8143d2fb;
  wire al_6f31a76;
  wire al_c5966d4f;
  wire al_e9ef2594;
  wire al_a7af1013;
  wire al_8d6e0488;
  wire al_4fc7a4fd;
  wire al_3660546c;
  wire al_cb807890;
  wire al_6d2e3f3;
  wire al_18c565c8;

  assign dBusAhb_HBURST[2] = 1'b0;
  assign dBusAhb_HBURST[1] = 1'b0;
  assign dBusAhb_HBURST[0] = 1'b0;
  assign dBusAhb_HPROT[3] = 1'b1;
  assign dBusAhb_HPROT[2] = 1'b1;
  assign dBusAhb_HPROT[1] = 1'b1;
  assign dBusAhb_HPROT[0] = 1'b1;
  assign dBusAhb_HSIZE[2] = 1'b0;
  assign dBusAhb_HSIZE[0] = al_bb6625de[1];
  assign dBusAhb_HTRANS[0] = 1'b0;
  assign iBusAhb_HADDR[31] = al_40185430[31];
  assign iBusAhb_HADDR[30] = al_40185430[30];
  assign iBusAhb_HADDR[29] = al_40185430[29];
  assign iBusAhb_HADDR[28] = al_40185430[28];
  assign iBusAhb_HADDR[27] = al_40185430[27];
  assign iBusAhb_HADDR[26] = al_40185430[26];
  assign iBusAhb_HADDR[25] = al_40185430[25];
  assign iBusAhb_HADDR[24] = al_40185430[24];
  assign iBusAhb_HADDR[23] = al_40185430[23];
  assign iBusAhb_HADDR[22] = al_40185430[22];
  assign iBusAhb_HADDR[21] = al_40185430[21];
  assign iBusAhb_HADDR[20] = al_40185430[20];
  assign iBusAhb_HADDR[19] = al_40185430[19];
  assign iBusAhb_HADDR[18] = al_40185430[18];
  assign iBusAhb_HADDR[17] = al_40185430[17];
  assign iBusAhb_HADDR[16] = al_40185430[16];
  assign iBusAhb_HADDR[15] = al_40185430[15];
  assign iBusAhb_HADDR[14] = al_40185430[14];
  assign iBusAhb_HADDR[13] = al_40185430[13];
  assign iBusAhb_HADDR[12] = al_40185430[12];
  assign iBusAhb_HADDR[11] = al_40185430[11];
  assign iBusAhb_HADDR[10] = al_40185430[10];
  assign iBusAhb_HADDR[9] = al_40185430[9];
  assign iBusAhb_HADDR[8] = al_40185430[8];
  assign iBusAhb_HADDR[7] = al_40185430[7];
  assign iBusAhb_HADDR[6] = al_40185430[6];
  assign iBusAhb_HADDR[5] = al_40185430[5];
  assign iBusAhb_HADDR[4] = al_40185430[4];
  assign iBusAhb_HADDR[3] = al_40185430[3];
  assign iBusAhb_HADDR[2] = al_40185430[2];
  assign iBusAhb_HADDR[1] = 1'b0;
  assign iBusAhb_HADDR[0] = 1'b0;
  assign iBusAhb_HBURST[2] = 1'b0;
  assign iBusAhb_HBURST[1] = 1'b0;
  assign iBusAhb_HBURST[0] = 1'b0;
  assign iBusAhb_HPROT[3] = 1'b1;
  assign iBusAhb_HPROT[2] = 1'b1;
  assign iBusAhb_HPROT[1] = 1'b1;
  assign iBusAhb_HPROT[0] = 1'b0;
  assign iBusAhb_HSIZE[2] = 1'b0;
  assign iBusAhb_HSIZE[1] = 1'b1;
  assign iBusAhb_HSIZE[0] = 1'b0;
  assign iBusAhb_HTRANS[1] = al_6897cc6d;
  assign iBusAhb_HTRANS[0] = 1'b0;
  assign iBusAhb_HWDATA[31] = 1'b0;
  assign iBusAhb_HWDATA[30] = 1'b0;
  assign iBusAhb_HWDATA[29] = 1'b0;
  assign iBusAhb_HWDATA[28] = 1'b0;
  assign iBusAhb_HWDATA[27] = 1'b0;
  assign iBusAhb_HWDATA[26] = 1'b0;
  assign iBusAhb_HWDATA[25] = 1'b0;
  assign iBusAhb_HWDATA[24] = 1'b0;
  assign iBusAhb_HWDATA[23] = 1'b0;
  assign iBusAhb_HWDATA[22] = 1'b0;
  assign iBusAhb_HWDATA[21] = 1'b0;
  assign iBusAhb_HWDATA[20] = 1'b0;
  assign iBusAhb_HWDATA[19] = 1'b0;
  assign iBusAhb_HWDATA[18] = 1'b0;
  assign iBusAhb_HWDATA[17] = 1'b0;
  assign iBusAhb_HWDATA[16] = 1'b0;
  assign iBusAhb_HWDATA[15] = 1'b0;
  assign iBusAhb_HWDATA[14] = 1'b0;
  assign iBusAhb_HWDATA[13] = 1'b0;
  assign iBusAhb_HWDATA[12] = 1'b0;
  assign iBusAhb_HWDATA[11] = 1'b0;
  assign iBusAhb_HWDATA[10] = 1'b0;
  assign iBusAhb_HWDATA[9] = 1'b0;
  assign iBusAhb_HWDATA[8] = 1'b0;
  assign iBusAhb_HWDATA[7] = 1'b0;
  assign iBusAhb_HWDATA[6] = 1'b0;
  assign iBusAhb_HWDATA[5] = 1'b0;
  assign iBusAhb_HWDATA[4] = 1'b0;
  assign iBusAhb_HWDATA[3] = 1'b0;
  assign iBusAhb_HWDATA[2] = 1'b0;
  assign iBusAhb_HWDATA[1] = 1'b0;
  assign iBusAhb_HWDATA[0] = 1'b0;
  assign iBusAhb_HWRITE = 1'b0;
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(E*~(F*~D*C*B)))"),
    .INIT(64'hffbfaaaaffffaaaa))
    al_56b6ffc1 (
    .a(INTERRUPT_i[0]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(al_d264c8ee[0]),
    .f(dBusAhb_HWDATA[0]),
    .o(al_f92bb470[0]));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(E*~(F*~D*C*B)))"),
    .INIT(64'hffbfaaaaffffaaaa))
    al_23e0ae21 (
    .a(INTERRUPT_i[1]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(al_d264c8ee[1]),
    .f(dBusAhb_HWDATA[1]),
    .o(al_f92bb470[1]));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(E*~(F*~D*C*B)))"),
    .INIT(64'hffbfaaaaffffaaaa))
    al_87804eb1 (
    .a(INTERRUPT_i[2]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(al_d264c8ee[2]),
    .f(dBusAhb_HWDATA[2]),
    .o(al_f92bb470[2]));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(E*~(F*~D*C*B)))"),
    .INIT(64'hffbfaaaaffffaaaa))
    al_ccaec426 (
    .a(INTERRUPT_i[3]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(al_d264c8ee[3]),
    .f(dBusAhb_HWDATA[3]),
    .o(al_f92bb470[3]));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(E*~(F*~D*C*B)))"),
    .INIT(64'hffbfaaaaffffaaaa))
    al_131276d0 (
    .a(INTERRUPT_i[4]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(al_d264c8ee[4]),
    .f(dBusAhb_HWDATA[4]),
    .o(al_f92bb470[4]));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(E*~(F*~D*C*B)))"),
    .INIT(64'hffbfaaaaffffaaaa))
    al_a8e6e1a8 (
    .a(INTERRUPT_i[5]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(al_d264c8ee[5]),
    .f(dBusAhb_HWDATA[5]),
    .o(al_f92bb470[5]));
  AL_DFF_X al_5d49c503 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f92bb470[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d264c8ee[0]));
  AL_DFF_X al_7a73169e (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f92bb470[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d264c8ee[1]));
  AL_DFF_X al_202a524 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f92bb470[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d264c8ee[2]));
  AL_DFF_X al_ac5a49ff (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f92bb470[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d264c8ee[3]));
  AL_DFF_X al_2950f550 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f92bb470[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d264c8ee[4]));
  AL_DFF_X al_ef9b17ec (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f92bb470[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d264c8ee[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_feffd2ed (
    .a(al_5d13c933[0]),
    .b(al_5d13c933[1]),
    .c(al_5d13c933[2]),
    .o(al_c0f2d5f7));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_837e34a8 (
    .a(al_921bc4ca),
    .b(al_831101f2[0]),
    .o(al_eb4cb082[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7aa33f0c (
    .a(al_921bc4ca),
    .b(al_831101f2[10]),
    .o(al_eb4cb082[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_8dbfc711 (
    .a(al_921bc4ca),
    .b(al_831101f2[11]),
    .o(al_eb4cb082[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_e3d0d98d (
    .a(al_921bc4ca),
    .b(al_831101f2[12]),
    .o(al_eb4cb082[12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_369f3e5b (
    .a(al_921bc4ca),
    .b(al_831101f2[13]),
    .o(al_eb4cb082[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_1ffb6bb3 (
    .a(al_921bc4ca),
    .b(al_831101f2[14]),
    .o(al_eb4cb082[14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_3f65f6ff (
    .a(al_921bc4ca),
    .b(al_831101f2[15]),
    .o(al_eb4cb082[15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_87391fe0 (
    .a(al_921bc4ca),
    .b(al_831101f2[16]),
    .o(al_eb4cb082[16]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_d3136c5e (
    .a(al_921bc4ca),
    .b(al_831101f2[17]),
    .o(al_eb4cb082[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_505819ff (
    .a(al_921bc4ca),
    .b(al_831101f2[18]),
    .o(al_eb4cb082[18]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_20b1ff5b (
    .a(al_921bc4ca),
    .b(al_831101f2[19]),
    .o(al_eb4cb082[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_90ad9e20 (
    .a(al_921bc4ca),
    .b(al_831101f2[1]),
    .o(al_eb4cb082[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_ace9e352 (
    .a(al_921bc4ca),
    .b(al_831101f2[20]),
    .o(al_eb4cb082[20]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_c7c85c75 (
    .a(al_921bc4ca),
    .b(al_831101f2[21]),
    .o(al_eb4cb082[21]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_2729c1ae (
    .a(al_921bc4ca),
    .b(al_831101f2[22]),
    .o(al_eb4cb082[22]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_58c1cc8 (
    .a(al_921bc4ca),
    .b(al_831101f2[23]),
    .o(al_eb4cb082[23]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_c01102ac (
    .a(al_921bc4ca),
    .b(al_831101f2[24]),
    .o(al_eb4cb082[24]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_541373a6 (
    .a(al_921bc4ca),
    .b(al_831101f2[25]),
    .o(al_eb4cb082[25]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_5b7695d6 (
    .a(al_921bc4ca),
    .b(al_831101f2[26]),
    .o(al_eb4cb082[26]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7ecc6313 (
    .a(al_921bc4ca),
    .b(al_831101f2[27]),
    .o(al_eb4cb082[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_f69f3429 (
    .a(al_ad9a3ca4[7]),
    .b(al_ad9a3ca4[22]),
    .c(al_ad9a3ca4[23]),
    .d(al_65949b4f[7]),
    .e(al_65949b4f[22]),
    .f(al_65949b4f[23]),
    .o(al_7ee9f8d));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_daf1f546 (
    .a(al_ad9a3ca4[2]),
    .b(al_ad9a3ca4[12]),
    .c(al_ad9a3ca4[13]),
    .d(al_65949b4f[2]),
    .e(al_65949b4f[12]),
    .f(al_65949b4f[13]),
    .o(al_942fb5b3));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_b60aba21 (
    .a(al_7ee9f8d),
    .b(al_bd909ea1),
    .c(al_80b19a9e),
    .d(al_be111ebc),
    .e(al_69da6feb),
    .f(al_942fb5b3),
    .o(al_31800d3e));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_6ba99054 (
    .a(al_ad9a3ca4[3]),
    .b(al_ad9a3ca4[17]),
    .c(al_ad9a3ca4[19]),
    .d(al_65949b4f[3]),
    .e(al_65949b4f[17]),
    .f(al_65949b4f[19]),
    .o(al_68c8085f));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_79833b91 (
    .a(al_ad9a3ca4[11]),
    .b(al_ad9a3ca4[14]),
    .c(al_ad9a3ca4[18]),
    .d(al_65949b4f[11]),
    .e(al_65949b4f[14]),
    .f(al_65949b4f[18]),
    .o(al_7a9d9124));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_6fa4432f (
    .a(al_ad9a3ca4[16]),
    .b(al_ad9a3ca4[25]),
    .c(al_ad9a3ca4[26]),
    .d(al_65949b4f[16]),
    .e(al_65949b4f[25]),
    .f(al_65949b4f[26]),
    .o(al_e85a2cb7));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_91b5b7a1 (
    .a(al_ad9a3ca4[4]),
    .b(al_ad9a3ca4[10]),
    .c(al_ad9a3ca4[21]),
    .d(al_65949b4f[4]),
    .e(al_65949b4f[10]),
    .f(al_65949b4f[21]),
    .o(al_ccef9e4c));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_efc57fd1 (
    .a(al_31800d3e),
    .b(al_68c8085f),
    .c(al_7a9d9124),
    .d(al_e85a2cb7),
    .e(al_ccef9e4c),
    .o(al_2e06c46d));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_9164e463 (
    .a(al_2e06c46d),
    .b(al_ad9a3ca4[30]),
    .o(al_921bc4ca));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_b8edd229 (
    .a(al_921bc4ca),
    .b(al_831101f2[28]),
    .o(al_eb4cb082[28]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_5600a9b1 (
    .a(al_ad9a3ca4[5]),
    .b(al_ad9a3ca4[6]),
    .c(al_ad9a3ca4[8]),
    .d(al_65949b4f[5]),
    .e(al_65949b4f[6]),
    .f(al_65949b4f[8]),
    .o(al_bd909ea1));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_78637da9 (
    .a(al_ad9a3ca4[15]),
    .b(al_ad9a3ca4[24]),
    .c(al_ad9a3ca4[29]),
    .d(al_65949b4f[15]),
    .e(al_65949b4f[24]),
    .f(al_65949b4f[29]),
    .o(al_80b19a9e));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_6dfa2f25 (
    .a(al_ad9a3ca4[0]),
    .b(al_ad9a3ca4[27]),
    .c(al_ad9a3ca4[28]),
    .d(al_65949b4f[0]),
    .e(al_65949b4f[27]),
    .f(al_65949b4f[28]),
    .o(al_be111ebc));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_6273388a (
    .a(al_ad9a3ca4[1]),
    .b(al_ad9a3ca4[9]),
    .c(al_ad9a3ca4[20]),
    .d(al_65949b4f[1]),
    .e(al_65949b4f[9]),
    .f(al_65949b4f[20]),
    .o(al_69da6feb));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_e1254103 (
    .a(al_921bc4ca),
    .b(al_831101f2[29]),
    .o(al_eb4cb082[29]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_78acc29d (
    .a(al_921bc4ca),
    .b(al_831101f2[2]),
    .o(al_eb4cb082[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_64225700 (
    .a(al_921bc4ca),
    .b(al_831101f2[3]),
    .o(al_eb4cb082[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_fd7271f0 (
    .a(al_921bc4ca),
    .b(al_831101f2[4]),
    .o(al_eb4cb082[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_ef091c68 (
    .a(al_921bc4ca),
    .b(al_831101f2[5]),
    .o(al_eb4cb082[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_b6c2920d (
    .a(al_921bc4ca),
    .b(al_831101f2[6]),
    .o(al_eb4cb082[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_922bf48 (
    .a(al_921bc4ca),
    .b(al_831101f2[7]),
    .o(al_eb4cb082[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_ddac12d2 (
    .a(al_921bc4ca),
    .b(al_831101f2[8]),
    .o(al_eb4cb082[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7c9ae259 (
    .a(al_921bc4ca),
    .b(al_831101f2[9]),
    .o(al_eb4cb082[9]));
  AL_DFF_X al_b76793d1 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ce484726),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92eee380));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E)*~((~D*~C*B))+A*E*~((~D*~C*B))+~(A)*E*(~D*~C*B)+A*E*(~D*~C*B))"),
    .INIT(32'haaaeaaa2))
    al_8c5a47c (
    .a(al_92eee380),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(dBusAhb_HWDATA[0]),
    .o(al_ce484726));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*~(E*~D*C))*~(B*A))"),
    .INIT(64'hff8fffff88888888))
    al_34749bd5 (
    .a(al_2e06c46d),
    .b(al_ad9a3ca4[30]),
    .c(al_5d13c933[0]),
    .d(al_5d13c933[1]),
    .e(al_5d13c933[2]),
    .f(al_384c501e),
    .o(al_747f0d5b));
  AL_DFF_X al_d84a40c4 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_747f0d5b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_384c501e));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_c447bb95 (
    .a(1'b0),
    .o({al_6a01eacd,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8343d5ff (
    .a(al_65949b4f[0]),
    .b(1'b1),
    .c(al_6a01eacd),
    .o({al_9ab3fa7e,al_831101f2[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cec55056 (
    .a(al_65949b4f[1]),
    .b(1'b0),
    .c(al_9ab3fa7e),
    .o({al_45a5e4cd,al_831101f2[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ff0030be (
    .a(al_65949b4f[2]),
    .b(1'b0),
    .c(al_45a5e4cd),
    .o({al_5fde6364,al_831101f2[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fd297d0b (
    .a(al_65949b4f[3]),
    .b(1'b0),
    .c(al_5fde6364),
    .o({al_98083b2a,al_831101f2[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1bb11246 (
    .a(al_65949b4f[4]),
    .b(1'b0),
    .c(al_98083b2a),
    .o({al_b935f70,al_831101f2[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d7d7480e (
    .a(al_65949b4f[5]),
    .b(1'b0),
    .c(al_b935f70),
    .o({al_72cf4613,al_831101f2[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fa410a31 (
    .a(al_65949b4f[6]),
    .b(1'b0),
    .c(al_72cf4613),
    .o({al_65e27d78,al_831101f2[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e2b6e66a (
    .a(al_65949b4f[7]),
    .b(1'b0),
    .c(al_65e27d78),
    .o({al_33785de1,al_831101f2[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1a7cb081 (
    .a(al_65949b4f[8]),
    .b(1'b0),
    .c(al_33785de1),
    .o({al_a50da65e,al_831101f2[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a99283fa (
    .a(al_65949b4f[9]),
    .b(1'b0),
    .c(al_a50da65e),
    .o({al_caba2fac,al_831101f2[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_158f2044 (
    .a(al_65949b4f[10]),
    .b(1'b0),
    .c(al_caba2fac),
    .o({al_82b381ff,al_831101f2[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c532ee78 (
    .a(al_65949b4f[11]),
    .b(1'b0),
    .c(al_82b381ff),
    .o({al_33365b48,al_831101f2[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b256fb16 (
    .a(al_65949b4f[12]),
    .b(1'b0),
    .c(al_33365b48),
    .o({al_c2fc5aeb,al_831101f2[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f23fe9de (
    .a(al_65949b4f[13]),
    .b(1'b0),
    .c(al_c2fc5aeb),
    .o({al_6ab36ff1,al_831101f2[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4c1bf607 (
    .a(al_65949b4f[14]),
    .b(1'b0),
    .c(al_6ab36ff1),
    .o({al_dd2f78da,al_831101f2[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5f057670 (
    .a(al_65949b4f[15]),
    .b(1'b0),
    .c(al_dd2f78da),
    .o({al_8179cfdf,al_831101f2[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_93ad47bc (
    .a(al_65949b4f[16]),
    .b(1'b0),
    .c(al_8179cfdf),
    .o({al_45cc89d,al_831101f2[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cd738ee3 (
    .a(al_65949b4f[17]),
    .b(1'b0),
    .c(al_45cc89d),
    .o({al_7568a715,al_831101f2[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1913eea3 (
    .a(al_65949b4f[18]),
    .b(1'b0),
    .c(al_7568a715),
    .o({al_4609cf3c,al_831101f2[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dc6c49cc (
    .a(al_65949b4f[19]),
    .b(1'b0),
    .c(al_4609cf3c),
    .o({al_e181a464,al_831101f2[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ff8d6eda (
    .a(al_65949b4f[20]),
    .b(1'b0),
    .c(al_e181a464),
    .o({al_b1593081,al_831101f2[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6bcf45d3 (
    .a(al_65949b4f[21]),
    .b(1'b0),
    .c(al_b1593081),
    .o({al_50a1040b,al_831101f2[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c97feaf3 (
    .a(al_65949b4f[22]),
    .b(1'b0),
    .c(al_50a1040b),
    .o({al_3e563e21,al_831101f2[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_224029ec (
    .a(al_65949b4f[23]),
    .b(1'b0),
    .c(al_3e563e21),
    .o({al_899000eb,al_831101f2[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_13ea81aa (
    .a(al_65949b4f[24]),
    .b(1'b0),
    .c(al_899000eb),
    .o({al_1c92cde,al_831101f2[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1a573a31 (
    .a(al_65949b4f[25]),
    .b(1'b0),
    .c(al_1c92cde),
    .o({al_e846ab0b,al_831101f2[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f798ccff (
    .a(al_65949b4f[26]),
    .b(1'b0),
    .c(al_e846ab0b),
    .o({al_78f1e056,al_831101f2[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f551ac7f (
    .a(al_65949b4f[27]),
    .b(1'b0),
    .c(al_78f1e056),
    .o({al_7704555,al_831101f2[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2695ecae (
    .a(al_65949b4f[28]),
    .b(1'b0),
    .c(al_7704555),
    .o({al_6a3d23ee,al_831101f2[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_aa8c73f1 (
    .a(al_65949b4f[29]),
    .b(1'b0),
    .c(al_6a3d23ee),
    .o({open_n3,al_831101f2[29]}));
  AL_DFF_X al_f7d0c35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[8]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[8]));
  AL_DFF_X al_785e84f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[9]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[9]));
  AL_DFF_X al_b8fb8ba5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[10]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[10]));
  AL_DFF_X al_a3368cef (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[11]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[11]));
  AL_DFF_X al_d73e99fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[12]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[12]));
  AL_DFF_X al_2449ecf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[13]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[13]));
  AL_DFF_X al_8b66cdea (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[14]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[14]));
  AL_DFF_X al_233deae9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[15]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[15]));
  AL_DFF_X al_b5d53eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[16]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[16]));
  AL_DFF_X al_362103c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[17]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[17]));
  AL_DFF_X al_460584bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[0]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[0]));
  AL_DFF_X al_6d89b5ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[18]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[18]));
  AL_DFF_X al_96585baf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[19]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[19]));
  AL_DFF_X al_2533ef4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[20]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[20]));
  AL_DFF_X al_4ed0fa49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[21]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[21]));
  AL_DFF_X al_e53f0ddf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[22]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[22]));
  AL_DFF_X al_10afa77e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[23]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[23]));
  AL_DFF_X al_1a348928 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[24]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[24]));
  AL_DFF_X al_6da0ad1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[25]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[25]));
  AL_DFF_X al_866dcc60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[26]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[26]));
  AL_DFF_X al_527c630a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[27]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[27]));
  AL_DFF_X al_145d0777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[1]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[1]));
  AL_DFF_X al_6485110b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[28]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[28]));
  AL_DFF_X al_bc557bad (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[29]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[29]));
  AL_DFF_X al_9b7f00cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cffac9df),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c5dfaf6[30]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_609308ad (
    .a(al_dc5ae5dc),
    .b(dBusAhb_HADDR[2]),
    .o(al_e84a0f1e));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_6f6e9f02 (
    .a(al_e84a0f1e),
    .b(al_ece70a8c),
    .c(al_ad9a3ca4[30]),
    .o(al_cffac9df));
  AL_DFF_X al_c4459ccd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[2]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[2]));
  AL_DFF_X al_5cfb2aaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[3]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[3]));
  AL_DFF_X al_ba9d086 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[4]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[4]));
  AL_DFF_X al_7219dadf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[5]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[5]));
  AL_DFF_X al_a6637fa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[6]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[6]));
  AL_DFF_X al_b0b52b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5d92ff7c[7]),
    .en(1'b1),
    .sr(~al_ece70a8c),
    .ss(1'b0),
    .q(al_7c5dfaf6[7]));
  AL_DFF_X al_e7d02df (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[8]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[8]));
  AL_DFF_X al_b7cf0b6a (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[9]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[9]));
  AL_DFF_X al_2262dc3f (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[10]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[10]));
  AL_DFF_X al_89a1b56b (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[11]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[11]));
  AL_DFF_X al_ebbbff5a (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[12]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[12]));
  AL_DFF_X al_cffeb3f4 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[13]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[13]));
  AL_DFF_X al_cffa3a38 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[14]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[14]));
  AL_DFF_X al_80a9b6b9 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[15]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[15]));
  AL_DFF_X al_5870fe1b (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[16]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[16]));
  AL_DFF_X al_508471e9 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[17]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[17]));
  AL_DFF_X al_125e7198 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[0]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[0]));
  AL_DFF_X al_7abcf8da (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[18]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[18]));
  AL_DFF_X al_112cb79e (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[19]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[19]));
  AL_DFF_X al_fa6bef54 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[20]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[20]));
  AL_DFF_X al_89994ba3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[21]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[21]));
  AL_DFF_X al_64dd9d42 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[22]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[22]));
  AL_DFF_X al_bcaca990 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[23]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[23]));
  AL_DFF_X al_8fd57143 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[24]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[24]));
  AL_DFF_X al_840fe4ad (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[25]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[25]));
  AL_DFF_X al_e176308c (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[26]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[26]));
  AL_DFF_X al_eec835da (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[27]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[27]));
  AL_DFF_X al_4d41a46e (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[1]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[1]));
  AL_DFF_X al_d67e6455 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[28]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[28]));
  AL_DFF_X al_41733a48 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[29]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[29]));
  AL_DFF_X al_3fbf66f3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[31]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[30]));
  AL_DFF_X al_274c614c (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[2]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[2]));
  AL_DFF_X al_981b99a9 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[3]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[3]));
  AL_DFF_X al_9c081c56 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[4]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[4]));
  AL_DFF_X al_da5e0833 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[5]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[5]));
  AL_DFF_X al_b1188847 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[6]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[6]));
  AL_DFF_X al_21486c2c (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(dBusAhb_HWDATA[7]),
    .en(al_c0f2d5f7),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad9a3ca4[7]));
  AL_DFF_X al_3c71b57c (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[8]));
  AL_DFF_X al_a1830718 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[9]));
  AL_DFF_X al_8395a509 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[10]));
  AL_DFF_X al_603bc786 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[11]));
  AL_DFF_X al_a270b6f7 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[12]));
  AL_DFF_X al_93b00bf2 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[13]));
  AL_DFF_X al_a3591445 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[14]));
  AL_DFF_X al_669f573d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[15]));
  AL_DFF_X al_dbe26d06 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[16]));
  AL_DFF_X al_7da73cf5 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[17]));
  AL_DFF_X al_8e758e5c (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[0]));
  AL_DFF_X al_72ec8310 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[18]));
  AL_DFF_X al_b1e5df84 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[19]));
  AL_DFF_X al_6baff0c4 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[20]));
  AL_DFF_X al_3ed917eb (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[21]));
  AL_DFF_X al_c709a462 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[22]));
  AL_DFF_X al_e6f0e013 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[23]));
  AL_DFF_X al_6206e91 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[24]));
  AL_DFF_X al_815d6252 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[25]));
  AL_DFF_X al_e6ff3674 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[26]));
  AL_DFF_X al_cb2af375 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[27]));
  AL_DFF_X al_a515cd44 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[1]));
  AL_DFF_X al_8507d07d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[28]));
  AL_DFF_X al_4ab09c3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[29]));
  AL_DFF_X al_82802507 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[2]));
  AL_DFF_X al_326fdba2 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[3]));
  AL_DFF_X al_1a91c1f6 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[4]));
  AL_DFF_X al_3a3fcaf2 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[5]));
  AL_DFF_X al_18ecf3fc (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[6]));
  AL_DFF_X al_76fc2664 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(TIM_CLK),
    .d(al_eb4cb082[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65949b4f[7]));
  AL_DFF_X al_1735245f (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_932f8140),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e108f0ff[0]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E)*~((~D*C*~B))+A*E*~((~D*C*~B))+~(A)*E*(~D*C*~B)+A*E*(~D*C*~B))"),
    .INIT(32'haabaaa8a))
    al_83c91e3c (
    .a(al_e108f0ff[5]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(dBusAhb_HWDATA[5]),
    .o(al_99e052bc));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E)*~((~D*C*~B))+A*E*~((~D*C*~B))+~(A)*E*(~D*C*~B)+A*E*(~D*C*~B))"),
    .INIT(32'haabaaa8a))
    al_41937136 (
    .a(al_e108f0ff[0]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(dBusAhb_HWDATA[0]),
    .o(al_932f8140));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E)*~((~D*C*~B))+A*E*~((~D*C*~B))+~(A)*E*(~D*C*~B)+A*E*(~D*C*~B))"),
    .INIT(32'haabaaa8a))
    al_2104e9d7 (
    .a(al_e108f0ff[1]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(dBusAhb_HWDATA[1]),
    .o(al_fa1d7661));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E)*~((~D*C*~B))+A*E*~((~D*C*~B))+~(A)*E*(~D*C*~B)+A*E*(~D*C*~B))"),
    .INIT(32'haabaaa8a))
    al_3eb3a892 (
    .a(al_e108f0ff[2]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(dBusAhb_HWDATA[2]),
    .o(al_6f8c3f2d));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E)*~((~D*C*~B))+A*E*~((~D*C*~B))+~(A)*E*(~D*C*~B)+A*E*(~D*C*~B))"),
    .INIT(32'haabaaa8a))
    al_362b5100 (
    .a(al_e108f0ff[3]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(dBusAhb_HWDATA[3]),
    .o(al_917164b4));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E)*~((~D*C*~B))+A*E*~((~D*C*~B))+~(A)*E*(~D*C*~B)+A*E*(~D*C*~B))"),
    .INIT(32'haabaaa8a))
    al_a268917e (
    .a(al_e108f0ff[4]),
    .b(al_5d13c933[0]),
    .c(al_5d13c933[1]),
    .d(al_5d13c933[2]),
    .e(dBusAhb_HWDATA[4]),
    .o(al_5ce11e05));
  AL_DFF_X al_ce134b28 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_fa1d7661),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e108f0ff[1]));
  AL_DFF_X al_df831760 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f8c3f2d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e108f0ff[2]));
  AL_DFF_X al_6e1ab3c9 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_917164b4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e108f0ff[3]));
  AL_DFF_X al_c2cac4c3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5ce11e05),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e108f0ff[4]));
  AL_DFF_X al_8311080d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_99e052bc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e108f0ff[5]));
  AL_DFF_X al_ec018347 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_24e92378[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d13c933[0]));
  AL_DFF_X al_fb271432 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_24e92378[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d13c933[1]));
  AL_DFF_X al_4dcac4e (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_24e92378[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d13c933[2]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_3bf48138 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[15]),
    .d(al_65949b4f[15]),
    .o(al_5d92ff7c[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_214a3ee2 (
    .a(al_63842eca),
    .b(dBusAhb_HADDR[14]),
    .c(dBusAhb_HADDR[13]),
    .o(al_8f7c15b2));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    al_5d09ac99 (
    .a(al_8f7c15b2),
    .b(dBusAhb_HADDR[2]),
    .c(al_e108f0ff[1]),
    .d(al_d264c8ee[1]),
    .o(al_133c9e7c));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(E*C)*~(D*A))"),
    .INIT(32'hfefceecc))
    al_e8d1ac69 (
    .a(al_e84a0f1e),
    .b(al_133c9e7c),
    .c(al_a7747a86),
    .d(al_ad9a3ca4[1]),
    .e(al_65949b4f[1]),
    .o(al_5d92ff7c[1]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    al_e9e4b783 (
    .a(al_8f7c15b2),
    .b(dBusAhb_HADDR[2]),
    .c(al_e108f0ff[2]),
    .d(al_d264c8ee[2]),
    .o(al_c71e5d62));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(E*C)*~(D*A))"),
    .INIT(32'hfefceecc))
    al_20bdb184 (
    .a(al_e84a0f1e),
    .b(al_c71e5d62),
    .c(al_a7747a86),
    .d(al_ad9a3ca4[2]),
    .e(al_65949b4f[2]),
    .o(al_5d92ff7c[2]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    al_beec1db4 (
    .a(al_8f7c15b2),
    .b(dBusAhb_HADDR[2]),
    .c(al_e108f0ff[3]),
    .d(al_d264c8ee[3]),
    .o(al_a2c0d252));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(E*C)*~(D*A))"),
    .INIT(32'hfefceecc))
    al_109e1ecc (
    .a(al_e84a0f1e),
    .b(al_a2c0d252),
    .c(al_a7747a86),
    .d(al_ad9a3ca4[3]),
    .e(al_65949b4f[3]),
    .o(al_5d92ff7c[3]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    al_3fad109c (
    .a(al_8f7c15b2),
    .b(dBusAhb_HADDR[2]),
    .c(al_e108f0ff[4]),
    .d(al_d264c8ee[4]),
    .o(al_9bc5b10b));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(E*C)*~(D*A))"),
    .INIT(32'hfefceecc))
    al_999d9e80 (
    .a(al_e84a0f1e),
    .b(al_9bc5b10b),
    .c(al_a7747a86),
    .d(al_ad9a3ca4[4]),
    .e(al_65949b4f[4]),
    .o(al_5d92ff7c[4]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    al_59aeb729 (
    .a(al_8f7c15b2),
    .b(dBusAhb_HADDR[2]),
    .c(al_e108f0ff[5]),
    .d(al_d264c8ee[5]),
    .o(al_1df2c985));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(E*C)*~(D*A))"),
    .INIT(32'hfefceecc))
    al_7b8b28a6 (
    .a(al_e84a0f1e),
    .b(al_1df2c985),
    .c(al_a7747a86),
    .d(al_ad9a3ca4[5]),
    .e(al_65949b4f[5]),
    .o(al_5d92ff7c[5]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_667810a2 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[6]),
    .d(al_65949b4f[6]),
    .o(al_5d92ff7c[6]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_580e1db9 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[7]),
    .d(al_65949b4f[7]),
    .o(al_5d92ff7c[7]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_f64c18e6 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[8]),
    .d(al_65949b4f[8]),
    .o(al_5d92ff7c[8]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_49f31dde (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[9]),
    .d(al_65949b4f[9]),
    .o(al_5d92ff7c[9]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_fd2febd8 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[10]),
    .d(al_65949b4f[10]),
    .o(al_5d92ff7c[10]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_2d06178c (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[11]),
    .d(al_65949b4f[11]),
    .o(al_5d92ff7c[11]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_38510224 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[12]),
    .d(al_65949b4f[12]),
    .o(al_5d92ff7c[12]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_5ebeb751 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[13]),
    .d(al_65949b4f[13]),
    .o(al_5d92ff7c[13]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_22a60f0e (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[14]),
    .d(al_65949b4f[14]),
    .o(al_5d92ff7c[14]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_66cd3402 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[16]),
    .d(al_65949b4f[16]),
    .o(al_5d92ff7c[16]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_eadba97b (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[17]),
    .d(al_65949b4f[17]),
    .o(al_5d92ff7c[17]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_76f3c45 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[18]),
    .d(al_65949b4f[18]),
    .o(al_5d92ff7c[18]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_9a942910 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[19]),
    .d(al_65949b4f[19]),
    .o(al_5d92ff7c[19]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_4cdf5fce (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[20]),
    .d(al_65949b4f[20]),
    .o(al_5d92ff7c[20]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_6dcdc857 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[21]),
    .d(al_65949b4f[21]),
    .o(al_5d92ff7c[21]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_632c430b (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[22]),
    .d(al_65949b4f[22]),
    .o(al_5d92ff7c[22]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_e5f69ece (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[23]),
    .d(al_65949b4f[23]),
    .o(al_5d92ff7c[23]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_a5b8174b (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[24]),
    .d(al_65949b4f[24]),
    .o(al_5d92ff7c[24]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_fd281677 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[25]),
    .d(al_65949b4f[25]),
    .o(al_5d92ff7c[25]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_43d238e8 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[26]),
    .d(al_65949b4f[26]),
    .o(al_5d92ff7c[26]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_cd4760e6 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[27]),
    .d(al_65949b4f[27]),
    .o(al_5d92ff7c[27]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_ed846854 (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[28]),
    .d(al_65949b4f[28]),
    .o(al_5d92ff7c[28]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    al_b8684c7e (
    .a(al_e84a0f1e),
    .b(al_a7747a86),
    .c(al_ad9a3ca4[29]),
    .d(al_65949b4f[29]),
    .o(al_5d92ff7c[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hcacbcecffafbfeff))
    al_a36f6be9 (
    .a(dBusAhb_HADDR[2]),
    .b(dBusAhb_HADDR[14]),
    .c(dBusAhb_HADDR[13]),
    .d(al_92eee380),
    .e(al_ad9a3ca4[0]),
    .f(al_e108f0ff[0]),
    .o(al_a99e75eb));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(~F*D)*~C*B)*~(E*A))"),
    .INIT(64'haeae0c0caaae000c))
    al_c5f97b8d (
    .a(al_a7747a86),
    .b(al_63842eca),
    .c(al_a99e75eb),
    .d(dBusAhb_HADDR[2]),
    .e(al_65949b4f[0]),
    .f(al_d264c8ee[0]),
    .o(al_5d92ff7c[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_312a7799 (
    .a(al_18077581[2]),
    .b(al_2cbb16b4[2]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(~B*~(C*(~(D)*~(E)*~(F)+D*E*~(F)+D*~(E)*F))))"),
    .INIT(64'h8888a888a88888a8))
    al_4a10f384 (
    .a(al_9c367b3e),
    .b(al_a7747a86),
    .c(al_63842eca),
    .d(dBusAhb_HADDR[2]),
    .e(dBusAhb_HADDR[14]),
    .f(dBusAhb_HADDR[13]),
    .o(al_24e92378[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_14a009f9 (
    .a(dBusAhb_HADDR[4]),
    .b(dBusAhb_HADDR[9]),
    .c(dBusAhb_HADDR[10]),
    .d(dBusAhb_HADDR[11]),
    .o(al_4aafd23e));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    al_e16a803a (
    .a(al_4aafd23e),
    .b(dBusAhb_HADDR[2]),
    .c(dBusAhb_HADDR[7]),
    .d(dBusAhb_HADDR[8]),
    .o(al_36b19484));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    al_a7aee661 (
    .a(dBusAhb_HADDR[15]),
    .b(dBusAhb_HADDR[14]),
    .c(dBusAhb_HADDR[13]),
    .d(dBusAhb_HADDR[12]),
    .o(al_3e310318));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_bc9a4143 (
    .a(al_36b19484),
    .b(al_3e310318),
    .c(dBusAhb_HADDR[3]),
    .d(dBusAhb_HADDR[5]),
    .e(dBusAhb_HADDR[6]),
    .o(al_a7747a86));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4c35b54d (
    .a(al_18077581[31]),
    .b(al_2cbb16b4[31]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_60b81e64 (
    .a(al_18077581[22]),
    .b(al_2cbb16b4[22]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e5ce824 (
    .a(al_18077581[21]),
    .b(al_2cbb16b4[21]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5cc5f92f (
    .a(al_18077581[20]),
    .b(al_2cbb16b4[20]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_922ae57a (
    .a(al_18077581[19]),
    .b(al_2cbb16b4[19]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9d95cedc (
    .a(al_18077581[18]),
    .b(al_2cbb16b4[18]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_99b67513 (
    .a(al_18077581[17]),
    .b(al_2cbb16b4[17]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_6fda9d31 (
    .a(al_18077581[16]),
    .b(al_2cbb16b4[16]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_97053d05 (
    .a(al_18077581[15]),
    .b(al_2cbb16b4[15]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_28ef160b (
    .a(al_18077581[14]),
    .b(al_2cbb16b4[14]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7e273412 (
    .a(al_18077581[13]),
    .b(al_2cbb16b4[13]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e2a78182 (
    .a(al_18077581[30]),
    .b(al_2cbb16b4[30]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_eb1399dd (
    .a(al_18077581[12]),
    .b(al_2cbb16b4[12]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1dd2bd24 (
    .a(al_18077581[4]),
    .b(al_2cbb16b4[4]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_80616e49 (
    .a(al_18077581[3]),
    .b(al_2cbb16b4[3]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_15816413 (
    .a(al_18077581[5]),
    .b(al_2cbb16b4[5]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_dda8388a (
    .a(al_18077581[6]),
    .b(al_2cbb16b4[6]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_236ce2b8 (
    .a(al_18077581[7]),
    .b(al_2cbb16b4[7]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2c992d5b (
    .a(al_18077581[8]),
    .b(al_2cbb16b4[8]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_739c18c8 (
    .a(al_18077581[9]),
    .b(al_2cbb16b4[9]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_9431e1d8 (
    .a(al_18077581[10]),
    .b(al_2cbb16b4[10]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1d8e2e5d (
    .a(al_18077581[11]),
    .b(al_2cbb16b4[11]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_de99cf39 (
    .a(al_18077581[29]),
    .b(al_2cbb16b4[29]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[29]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_778d9d52 (
    .a(dBusAhb_HADDR[27]),
    .b(dBusAhb_HADDR[26]),
    .c(dBusAhb_HADDR[25]),
    .d(dBusAhb_HADDR[24]),
    .e(dBusAhb_HADDR[23]),
    .f(dBusAhb_HADDR[22]),
    .o(al_2fcd16aa));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_580703d7 (
    .a(dBusAhb_HADDR[19]),
    .b(dBusAhb_HADDR[18]),
    .c(dBusAhb_HADDR[17]),
    .d(dBusAhb_HADDR[16]),
    .o(al_82aaac97));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_51387259 (
    .a(dBusAhb_HADDR[31]),
    .b(dBusAhb_HADDR[30]),
    .c(dBusAhb_HADDR[29]),
    .d(dBusAhb_HADDR[28]),
    .o(al_dca31e55));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_b83461d2 (
    .a(al_2fcd16aa),
    .b(al_82aaac97),
    .c(al_dca31e55),
    .d(dBusAhb_HADDR[21]),
    .e(dBusAhb_HADDR[20]),
    .o(al_ece70a8c));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_7c29fff2 (
    .a(dBusAhb_HADDR[3]),
    .b(dBusAhb_HADDR[9]),
    .c(dBusAhb_HADDR[10]),
    .d(dBusAhb_HADDR[11]),
    .o(al_1cf6c96));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_d621a8b0 (
    .a(dBusAhb_HADDR[15]),
    .b(dBusAhb_HADDR[12]),
    .c(dBusAhb_HADDR[5]),
    .d(dBusAhb_HADDR[6]),
    .o(al_a4a54bdd));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_79d61ebf (
    .a(al_18077581[28]),
    .b(al_2cbb16b4[28]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[28]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_9e19722d (
    .a(al_1cf6c96),
    .b(al_a4a54bdd),
    .c(dBusAhb_HADDR[4]),
    .d(dBusAhb_HADDR[7]),
    .e(dBusAhb_HADDR[8]),
    .o(al_63842eca));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*~C*~B*~A)"),
    .INIT(64'h0100000000000000))
    al_cecf17b8 (
    .a(al_7bc36116),
    .b(al_bec39e4d),
    .c(al_6ec8afa5),
    .d(al_c572d1c7),
    .e(al_32fedef4),
    .f(al_523cde28),
    .o(al_1a09507b));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_db9f5d90 (
    .a(al_ece70a8c),
    .b(al_1a09507b),
    .c(dBusAhb_HWRITE),
    .o(al_9c367b3e));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    al_6d8ac461 (
    .a(al_9c367b3e),
    .b(al_63842eca),
    .c(dBusAhb_HADDR[14]),
    .d(dBusAhb_HADDR[13]),
    .o(al_24e92378[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_fb166b22 (
    .a(al_18077581[27]),
    .b(al_2cbb16b4[27]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_39776367 (
    .a(al_18077581[26]),
    .b(al_2cbb16b4[26]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_71b9ff42 (
    .a(al_18077581[25]),
    .b(al_2cbb16b4[25]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_99d2a72a (
    .a(al_18077581[24]),
    .b(al_2cbb16b4[24]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_61f17297 (
    .a(al_18077581[23]),
    .b(al_2cbb16b4[23]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[23]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_92d59d30 (
    .a(al_63842eca),
    .b(dBusAhb_HADDR[14]),
    .c(dBusAhb_HADDR[13]),
    .o(al_dc5ae5dc));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    al_f7704315 (
    .a(al_9c367b3e),
    .b(al_dc5ae5dc),
    .c(al_a7747a86),
    .o(al_24e92378[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_49ae92d8 (
    .a(al_a3a8b68d),
    .b(al_85a2bdb0[0]),
    .o(al_4d9a3d8e[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf7b3d591e6a2c480))
    al_63ab7b7b (
    .a(al_289dceb2),
    .b(al_dc412458),
    .c(al_4d9a3d8e[0]),
    .d(al_45e5d9f7[0]),
    .e(al_e03b3126[0]),
    .f(al_bfc96350[0]),
    .o(al_3dcca8e[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_e9e8e285 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[10]),
    .d(al_126b3afd[10]),
    .e(al_85a2bdb0[10]),
    .f(al_e03b3126[10]),
    .o(al_b1924903));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_8a4b4d53 (
    .a(al_b1924903),
    .b(al_6ec8afa5),
    .c(al_bfc96350[10]),
    .o(al_3dcca8e[10]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_fd19e711 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[11]),
    .d(al_126b3afd[11]),
    .e(al_85a2bdb0[11]),
    .o(al_569f263c));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_2aca5285 (
    .a(al_569f263c),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[11]),
    .e(al_bfc96350[11]),
    .o(al_3dcca8e[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_f058eee2 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[12]),
    .d(al_126b3afd[12]),
    .e(al_85a2bdb0[12]),
    .f(al_bb6625de[1]),
    .o(al_36303862));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_8ba6918f (
    .a(al_36303862),
    .b(al_6ec8afa5),
    .c(al_bfc96350[12]),
    .o(al_3dcca8e[12]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_d0600fb4 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[13]),
    .d(al_126b3afd[13]),
    .e(al_85a2bdb0[13]),
    .o(al_bc831201));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_75ae133a (
    .a(al_bc831201),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(dBusAhb_HSIZE[1]),
    .e(al_bfc96350[13]),
    .o(al_3dcca8e[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_83c8989f (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[14]),
    .d(al_126b3afd[14]),
    .e(al_85a2bdb0[14]),
    .f(al_e03b3126[14]),
    .o(al_1b5c5256));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_21d70052 (
    .a(al_1b5c5256),
    .b(al_6ec8afa5),
    .c(al_bfc96350[14]),
    .o(al_3dcca8e[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_3d1a96f6 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[15]),
    .d(al_126b3afd[15]),
    .e(al_85a2bdb0[15]),
    .f(al_e03b3126[15]),
    .o(al_9ce6f9ae));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_a3b356d7 (
    .a(al_9ce6f9ae),
    .b(al_6ec8afa5),
    .c(al_bfc96350[15]),
    .o(al_3dcca8e[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_240dac4b (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[16]),
    .d(al_126b3afd[16]),
    .e(al_85a2bdb0[16]),
    .o(al_d66e22dd));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_e5ebd314 (
    .a(al_d66e22dd),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[16]),
    .e(al_bfc96350[16]),
    .o(al_3dcca8e[16]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_b0071850 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[17]),
    .d(al_126b3afd[17]),
    .e(al_85a2bdb0[17]),
    .o(al_278217fa));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_1486e6e1 (
    .a(al_278217fa),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[17]),
    .e(al_bfc96350[17]),
    .o(al_3dcca8e[17]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_1dbcd071 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[18]),
    .d(al_126b3afd[18]),
    .e(al_85a2bdb0[18]),
    .o(al_f8b84ed9));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_18d0d739 (
    .a(al_f8b84ed9),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[18]),
    .e(al_bfc96350[18]),
    .o(al_3dcca8e[18]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_db58a61 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[19]),
    .d(al_126b3afd[19]),
    .e(al_85a2bdb0[19]),
    .f(al_e03b3126[19]),
    .o(al_b6d6e907));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_87d64234 (
    .a(al_b6d6e907),
    .b(al_6ec8afa5),
    .c(al_bfc96350[19]),
    .o(al_3dcca8e[19]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    al_993885f2 (
    .a(al_a8151162),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .o(al_289dceb2));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_842e604f (
    .a(al_6ec8afa5),
    .b(al_a5849610),
    .o(al_dc412458));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_72e5f0ab (
    .a(al_a3a8b68d),
    .b(al_85a2bdb0[1]),
    .o(al_4d9a3d8e[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf7b3d591e6a2c480))
    al_f40da571 (
    .a(al_289dceb2),
    .b(al_dc412458),
    .c(al_4d9a3d8e[1]),
    .d(al_45e5d9f7[1]),
    .e(al_e03b3126[1]),
    .f(al_bfc96350[1]),
    .o(al_3dcca8e[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_4e4f2697 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[20]),
    .d(al_126b3afd[20]),
    .e(al_85a2bdb0[20]),
    .o(al_44ee9376));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_4801d19a (
    .a(al_44ee9376),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[20]),
    .e(al_bfc96350[20]),
    .o(al_3dcca8e[20]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_c9d074f4 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[21]),
    .d(al_126b3afd[21]),
    .e(al_85a2bdb0[21]),
    .o(al_79fcc7dd));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_87e1b406 (
    .a(al_79fcc7dd),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[21]),
    .e(al_bfc96350[21]),
    .o(al_3dcca8e[21]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_5a5f0b73 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[22]),
    .d(al_126b3afd[22]),
    .e(al_85a2bdb0[22]),
    .o(al_f465aa2));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_123b074a (
    .a(al_f465aa2),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[22]),
    .e(al_bfc96350[22]),
    .o(al_3dcca8e[22]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_7bc20711 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[23]),
    .d(al_126b3afd[23]),
    .e(al_85a2bdb0[23]),
    .f(al_e03b3126[23]),
    .o(al_8675b08));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_4e9d2c1f (
    .a(al_8675b08),
    .b(al_6ec8afa5),
    .c(al_bfc96350[23]),
    .o(al_3dcca8e[23]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_4601a824 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[24]),
    .d(al_126b3afd[24]),
    .e(al_85a2bdb0[24]),
    .o(al_1e27127a));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_9ce742fa (
    .a(al_1e27127a),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[24]),
    .e(al_bfc96350[24]),
    .o(al_3dcca8e[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_b3a0f577 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[25]),
    .d(al_126b3afd[25]),
    .e(al_85a2bdb0[25]),
    .f(al_e03b3126[25]),
    .o(al_86608ce5));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_e00332c1 (
    .a(al_86608ce5),
    .b(al_6ec8afa5),
    .c(al_bfc96350[25]),
    .o(al_3dcca8e[25]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_280bc3da (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[26]),
    .d(al_126b3afd[26]),
    .e(al_85a2bdb0[26]),
    .o(al_dc741944));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_ca34f9d7 (
    .a(al_dc741944),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[26]),
    .e(al_bfc96350[26]),
    .o(al_3dcca8e[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_86181f62 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[27]),
    .d(al_126b3afd[27]),
    .e(al_85a2bdb0[27]),
    .f(al_e03b3126[27]),
    .o(al_730b0315));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_3f0569ca (
    .a(al_730b0315),
    .b(al_6ec8afa5),
    .c(al_bfc96350[27]),
    .o(al_3dcca8e[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_4b7abd95 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[28]),
    .d(al_126b3afd[28]),
    .e(al_85a2bdb0[28]),
    .f(al_e03b3126[28]),
    .o(al_14651309));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_5a6c7e08 (
    .a(al_14651309),
    .b(al_6ec8afa5),
    .c(al_bfc96350[28]),
    .o(al_3dcca8e[28]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b6e323d0 (
    .a(al_a8151162),
    .b(al_a5849610),
    .o(al_ce0d355f));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    al_f83bd9d0 (
    .a(al_a8151162),
    .b(al_a5849610),
    .c(al_a3a8b68d),
    .o(al_bd56460d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_ca996c9d (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[29]),
    .d(al_126b3afd[29]),
    .e(al_85a2bdb0[29]),
    .f(al_e03b3126[29]),
    .o(al_c0406dbc));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_d9991f4 (
    .a(al_c0406dbc),
    .b(al_6ec8afa5),
    .c(al_bfc96350[29]),
    .o(al_3dcca8e[29]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_3829a863 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[2]),
    .d(al_126b3afd[2]),
    .e(al_85a2bdb0[2]),
    .o(al_50c53403));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_f04e3a9f (
    .a(al_50c53403),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[2]),
    .e(al_bfc96350[2]),
    .o(al_3dcca8e[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_640e2688 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[30]),
    .d(al_126b3afd[30]),
    .e(al_85a2bdb0[30]),
    .o(al_36d679eb));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_5b32cfc1 (
    .a(al_36d679eb),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[30]),
    .e(al_bfc96350[30]),
    .o(al_3dcca8e[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_b884982a (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[31]),
    .d(al_126b3afd[31]),
    .e(al_85a2bdb0[31]),
    .f(al_e03b3126[31]),
    .o(al_e5ffe4ff));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_e6076f1c (
    .a(al_e5ffe4ff),
    .b(al_6ec8afa5),
    .c(al_bfc96350[31]),
    .o(al_3dcca8e[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_35085de4 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[3]),
    .d(al_126b3afd[3]),
    .e(al_85a2bdb0[3]),
    .f(al_e03b3126[3]),
    .o(al_f2fcadd6));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_9ccd85fd (
    .a(al_f2fcadd6),
    .b(al_6ec8afa5),
    .c(al_bfc96350[3]),
    .o(al_3dcca8e[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_9a93a783 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[4]),
    .d(al_126b3afd[4]),
    .e(al_85a2bdb0[4]),
    .f(al_e03b3126[4]),
    .o(al_7b2239bb));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_c079a1e6 (
    .a(al_7b2239bb),
    .b(al_6ec8afa5),
    .c(al_bfc96350[4]),
    .o(al_3dcca8e[4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_f389045a (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[5]),
    .d(al_126b3afd[5]),
    .e(al_85a2bdb0[5]),
    .o(al_c78a6044));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_3eab870c (
    .a(al_c78a6044),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(dBusAhb_HWRITE),
    .e(al_bfc96350[5]),
    .o(al_3dcca8e[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_85f4b77c (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[6]),
    .d(al_126b3afd[6]),
    .e(al_85a2bdb0[6]),
    .f(al_e03b3126[6]),
    .o(al_3cd3f418));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_a5f31d63 (
    .a(al_3cd3f418),
    .b(al_6ec8afa5),
    .c(al_bfc96350[6]),
    .o(al_3dcca8e[6]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_e0c93c4c (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[7]),
    .d(al_126b3afd[7]),
    .e(al_85a2bdb0[7]),
    .o(al_5c3a44f0));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_b018527f (
    .a(al_5c3a44f0),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[7]),
    .e(al_bfc96350[7]),
    .o(al_3dcca8e[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h048c26ae159d37bf))
    al_779aa076 (
    .a(al_ce0d355f),
    .b(al_bd56460d),
    .c(al_45e5d9f7[8]),
    .d(al_126b3afd[8]),
    .e(al_85a2bdb0[8]),
    .f(al_e03b3126[8]),
    .o(al_b5b0f369));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_c5d4ea38 (
    .a(al_b5b0f369),
    .b(al_6ec8afa5),
    .c(al_bfc96350[8]),
    .o(al_3dcca8e[8]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h024e135f))
    al_bbc06643 (
    .a(al_a8151162),
    .b(al_a3a8b68d),
    .c(al_45e5d9f7[9]),
    .d(al_126b3afd[9]),
    .e(al_85a2bdb0[9]),
    .o(al_41adb443));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*~(E)*~(B)+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*~(B)+~(~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))*E*B+~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C)*E*B)"),
    .INIT(32'hdfdc1310))
    al_75587900 (
    .a(al_41adb443),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e03b3126[9]),
    .e(al_bfc96350[9]),
    .o(al_3dcca8e[9]));
  AL_MAP_LUT6 #(
    .EQN("(~E*~B*~(C*~(~D*~(F*A))))"),
    .INIT(64'h0000031300000333))
    al_4d73b76 (
    .a(al_a8151162),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_a3a8b68d),
    .e(al_c85db05d),
    .f(al_7b80e496[0]),
    .o(al_319b4c4c));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    al_dba6d786 (
    .a(al_319b4c4c),
    .b(al_673a4598),
    .c(al_e3edcf1a),
    .d(al_501dbbdf),
    .o(al_9d1d880c[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(~D*A)))"),
    .INIT(16'hc0c8))
    al_bd3250f9 (
    .a(al_a8151162),
    .b(al_a5849610),
    .c(al_a3a8b68d),
    .d(al_7b80e496[1]),
    .o(al_f0561e92));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_b156a580 (
    .a(al_f0561e92),
    .b(al_6ec8afa5),
    .c(al_587b9831),
    .o(al_9d1d880c[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_d5336759 (
    .a(al_66ffb9),
    .b(al_a7b01c14[2]),
    .o(al_5fe8f9ad));
  AL_DFF_X al_b60b4fb0 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5fe8f9ad),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d2c853e));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*A))*~(C)+B*(D*A)*~(C)+~(B)*(D*A)*C+B*(D*A)*C)"),
    .INIT(16'hac0c))
    al_3f6f4207 (
    .a(al_66ffb9),
    .b(al_119831c0),
    .c(al_5a744f0f),
    .d(al_6f08d701),
    .o(al_9a3c3a5));
  AL_DFF_X al_daa7db0c (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9a3c3a5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b469f7cc));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(~F*~E)*~D*C)*~(B*A))"),
    .INIT(64'h88f888f888f88888))
    al_303b7292 (
    .a(al_119831c0),
    .b(al_5a744f0f),
    .c(al_9d63e9cd),
    .d(al_bb0cd305),
    .e(al_6ec8afa5),
    .f(al_d508bbc9),
    .o(al_d79e66b7));
  AL_DFF_X al_d05bbc48 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d79e66b7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d508bbc9));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    al_b3b23a73 (
    .a(al_9d63e9cd),
    .b(al_bb0cd305),
    .c(al_6ec8afa5),
    .d(al_d508bbc9),
    .o(al_5e3d90d7));
  AL_DFF_X al_fc6d9277 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5e3d90d7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6499e5fd));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_fd2a6515 (
    .a(al_6499e5fd),
    .b(al_8c0460e8),
    .o(al_c4074784));
  AL_DFF_X al_81a1220d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c4074784),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e275e81));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    al_9d422d25 (
    .a(al_da7f07ab),
    .b(al_aa37cfdb),
    .c(al_8869249d),
    .d(al_3697c94f),
    .o(al_89ab45b5));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    al_b2318e (
    .a(al_89ab45b5),
    .b(al_172eec6a),
    .c(al_a1a600b6),
    .o(al_4d82afcf));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(~C*A))"),
    .INIT(16'h3100))
    al_7d6e2cfd (
    .a(al_bec39e4d),
    .b(al_4d82afcf),
    .c(al_5e275e81),
    .d(al_ac1a4f11),
    .o(al_c871f2ad));
  AL_DFF_X al_b9d4d0eb (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c871f2ad),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b567677b));
  AL_DFF_X al_ce1624d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_4c590039),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ee8b2558));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    al_4564627c (
    .a(al_bec39e4d),
    .b(al_5e275e81),
    .c(al_ee8b2558),
    .o(al_4c590039));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(D*B)*~(E*A))"),
    .INIT(64'h0105030f115533ff))
    al_84b04f32 (
    .a(al_be8ea5e1),
    .b(al_4cc0b8dd),
    .c(al_7610b7fc),
    .d(al_1a8c7c22[0]),
    .e(al_ccabc055[0]),
    .f(al_97943858[0]),
    .o(al_193dedee));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    al_2fa1abaa (
    .a(al_193dedee),
    .b(al_235de557),
    .c(al_d19b9f6b),
    .d(al_41e76523[0]),
    .o(al_c0855656));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_e5a192ab (
    .a(al_c0855656),
    .b(al_18077581[0]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[0]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_a7a58c7b (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[0]),
    .c(al_c91705db),
    .d(al_ccabc055[0]),
    .e(al_e45b51d9[0]),
    .o(al_c28c3a52[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_f646befe (
    .a(al_555b0990[0]),
    .b(al_555b0990[1]),
    .c(al_407c8ac1),
    .o(al_18077581[10]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_3be6497 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[8]),
    .e(al_ccabc055[10]),
    .f(al_97943858[10]),
    .o(al_354f5999));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_36f3a5a9 (
    .a(al_354f5999),
    .b(al_18077581[10]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_cbb0a84b (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[10]),
    .d(al_ccabc055[10]),
    .e(al_e45b51d9[10]),
    .o(al_c28c3a52[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_2981ab2e (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[11]),
    .c(al_c91705db),
    .d(al_ccabc055[11]),
    .e(al_e45b51d9[11]),
    .o(al_c28c3a52[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_2613664b (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[12]),
    .c(al_c91705db),
    .d(al_ccabc055[12]),
    .e(al_e45b51d9[12]),
    .o(al_c28c3a52[12]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_aebae713 (
    .a(dBusAhb_HSIZE[1]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_c8ba6c61),
    .o(al_18077581[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_3985e72b (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[11]),
    .e(al_ccabc055[13]),
    .f(al_97943858[13]),
    .o(al_5914a559));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_ee7cce38 (
    .a(al_5914a559),
    .b(al_235de557),
    .o(al_85bef49));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_900f8552 (
    .a(al_85bef49),
    .b(al_18077581[13]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[13]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_593378c7 (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[13]),
    .c(al_c91705db),
    .d(al_ccabc055[13]),
    .e(al_e45b51d9[13]),
    .o(al_c28c3a52[13]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_76e8ebaf (
    .a(al_e03b3126[14]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_59be2ab1),
    .o(al_18077581[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_3e4aafdc (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[12]),
    .e(al_ccabc055[14]),
    .f(al_97943858[14]),
    .o(al_f6c8a5f0));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_b512d86a (
    .a(al_f6c8a5f0),
    .b(al_235de557),
    .o(al_94f9539));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_947dda89 (
    .a(al_94f9539),
    .b(al_18077581[14]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_d44bada0 (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[14]),
    .c(al_c91705db),
    .d(al_ccabc055[14]),
    .e(al_e45b51d9[14]),
    .o(al_c28c3a52[14]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_a20580f1 (
    .a(al_e03b3126[15]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_8488923),
    .o(al_18077581[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_b76ef0c9 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[13]),
    .e(al_ccabc055[15]),
    .f(al_97943858[15]),
    .o(al_f49386));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_b0fa0efb (
    .a(al_f49386),
    .b(al_18077581[15]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_768c2a0b (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[15]),
    .d(al_ccabc055[15]),
    .e(al_e45b51d9[15]),
    .o(al_c28c3a52[15]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_de22f88 (
    .a(al_e03b3126[16]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_5727b773),
    .o(al_18077581[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_33ea081c (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[14]),
    .e(al_ccabc055[16]),
    .f(al_97943858[16]),
    .o(al_bf987e25));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5f8dc364 (
    .a(al_bf987e25),
    .b(al_235de557),
    .o(al_b44f8827));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_3a205f21 (
    .a(al_b44f8827),
    .b(al_18077581[16]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[16]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_84f48336 (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[16]),
    .c(al_c91705db),
    .d(al_ccabc055[16]),
    .e(al_e45b51d9[16]),
    .o(al_c28c3a52[16]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_68444bc3 (
    .a(al_e03b3126[17]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_eead7739),
    .o(al_18077581[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_5be52a73 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[15]),
    .e(al_ccabc055[17]),
    .f(al_97943858[17]),
    .o(al_daaf28b4));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_2ff7dd3b (
    .a(al_daaf28b4),
    .b(al_18077581[17]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[17]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_6911867 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[17]),
    .d(al_ccabc055[17]),
    .e(al_e45b51d9[17]),
    .o(al_c28c3a52[17]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_e6cbea81 (
    .a(al_e03b3126[18]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_f430a5aa),
    .o(al_18077581[18]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_406a40ac (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[16]),
    .e(al_ccabc055[18]),
    .f(al_97943858[18]),
    .o(al_5c0f2717));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_fdc06a16 (
    .a(al_5c0f2717),
    .b(al_18077581[18]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[18]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_e8efecb8 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[18]),
    .d(al_ccabc055[18]),
    .e(al_e45b51d9[18]),
    .o(al_c28c3a52[18]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_951fbfb5 (
    .a(al_e03b3126[19]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_cd498e9f),
    .o(al_18077581[19]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_21122dc8 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[17]),
    .e(al_ccabc055[19]),
    .f(al_97943858[19]),
    .o(al_8a79ceb4));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_447d0845 (
    .a(al_8a79ceb4),
    .b(al_18077581[19]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[19]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_84a02c60 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[19]),
    .d(al_ccabc055[19]),
    .e(al_e45b51d9[19]),
    .o(al_c28c3a52[19]));
  AL_MAP_LUT6 #(
    .EQN("(~B*~A*~(F*D)*~(E*C))"),
    .INIT(64'h0001001101011111))
    al_aa769fdf (
    .a(al_235de557),
    .b(al_9c55c5c3),
    .c(al_d19b9f6b),
    .d(al_be8ea5e1),
    .e(al_41e76523[1]),
    .f(al_ccabc055[1]),
    .o(al_bdfc704c));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    al_5676c480 (
    .a(al_bdfc704c),
    .b(al_4cc0b8dd),
    .c(al_7610b7fc),
    .d(al_1a8c7c22[1]),
    .e(al_97943858[1]),
    .o(al_f4418953));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_f6245c6c (
    .a(al_f4418953),
    .b(al_18077581[1]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_fbaf7126 (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[1]),
    .c(al_c91705db),
    .d(al_ccabc055[1]),
    .e(al_e45b51d9[1]),
    .o(al_c28c3a52[1]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_75c5216 (
    .a(al_e03b3126[20]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_3656d228),
    .o(al_18077581[20]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_4dfabda4 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[18]),
    .e(al_ccabc055[20]),
    .f(al_97943858[20]),
    .o(al_65a874f0));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_4029dcde (
    .a(al_65a874f0),
    .b(al_18077581[20]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[20]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_353a5da9 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[20]),
    .d(al_ccabc055[20]),
    .e(al_e45b51d9[20]),
    .o(al_c28c3a52[20]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_5a1f14af (
    .a(al_e03b3126[21]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_30f08f9c),
    .o(al_18077581[21]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_6a8b5de3 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[19]),
    .e(al_ccabc055[21]),
    .f(al_97943858[21]),
    .o(al_80b925b7));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_6d5736bf (
    .a(al_80b925b7),
    .b(al_18077581[21]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[21]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_87e980e2 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[21]),
    .d(al_ccabc055[21]),
    .e(al_e45b51d9[21]),
    .o(al_c28c3a52[21]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_39bd823f (
    .a(al_e03b3126[22]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_bf6a3977),
    .o(al_18077581[22]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_960222f3 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[20]),
    .e(al_ccabc055[22]),
    .f(al_97943858[22]),
    .o(al_dfe3b0a5));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_72894401 (
    .a(al_dfe3b0a5),
    .b(al_235de557),
    .o(al_cb828215));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_18d30289 (
    .a(al_cb828215),
    .b(al_18077581[22]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[22]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_e7ea5737 (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[22]),
    .c(al_c91705db),
    .d(al_ccabc055[22]),
    .e(al_e45b51d9[22]),
    .o(al_c28c3a52[22]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_3c4a8115 (
    .a(al_e03b3126[23]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_2ede456b),
    .o(al_18077581[23]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_cc982075 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[21]),
    .e(al_ccabc055[23]),
    .f(al_97943858[23]),
    .o(al_ce80e68f));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_2d84471b (
    .a(al_ce80e68f),
    .b(al_18077581[23]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[23]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_d61d4ae3 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[23]),
    .d(al_ccabc055[23]),
    .e(al_e45b51d9[23]),
    .o(al_c28c3a52[23]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_a8404fc (
    .a(al_e03b3126[24]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_3a7c5a5),
    .o(al_18077581[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_e55155a9 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[22]),
    .e(al_ccabc055[24]),
    .f(al_97943858[24]),
    .o(al_14816c03));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_101e5f5a (
    .a(al_14816c03),
    .b(al_18077581[24]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[24]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_518b356d (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[24]),
    .d(al_ccabc055[24]),
    .e(al_e45b51d9[24]),
    .o(al_c28c3a52[24]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_65b06768 (
    .a(al_e03b3126[25]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_9b707062),
    .o(al_18077581[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_834ea514 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[23]),
    .e(al_ccabc055[25]),
    .f(al_97943858[25]),
    .o(al_6d174013));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_c9ab464b (
    .a(al_6d174013),
    .b(al_18077581[25]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[25]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_2fd2d86a (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[25]),
    .d(al_ccabc055[25]),
    .e(al_e45b51d9[25]),
    .o(al_c28c3a52[25]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_8e9d74f9 (
    .a(al_e03b3126[26]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_a69cec28),
    .o(al_18077581[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_fb81efb5 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[24]),
    .e(al_ccabc055[26]),
    .f(al_97943858[26]),
    .o(al_385f14));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_7f0b67a0 (
    .a(al_385f14),
    .b(al_235de557),
    .o(al_bb4f8966));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_b653a17f (
    .a(al_bb4f8966),
    .b(al_18077581[26]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[26]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_68178a1b (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[26]),
    .c(al_c91705db),
    .d(al_ccabc055[26]),
    .e(al_e45b51d9[26]),
    .o(al_c28c3a52[26]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_8cae4cc4 (
    .a(al_e03b3126[27]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_d78f6bd4),
    .o(al_18077581[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_484717d1 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[25]),
    .e(al_ccabc055[27]),
    .f(al_97943858[27]),
    .o(al_70fea121));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_a6d108ac (
    .a(al_70fea121),
    .b(al_18077581[27]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[27]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_faca0e17 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[27]),
    .d(al_ccabc055[27]),
    .e(al_e45b51d9[27]),
    .o(al_c28c3a52[27]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_b15beb4f (
    .a(al_e03b3126[28]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_cae21d2e),
    .o(al_18077581[28]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_1affd539 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[26]),
    .e(al_ccabc055[28]),
    .f(al_97943858[28]),
    .o(al_7750a3cd));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_83765894 (
    .a(al_7750a3cd),
    .b(al_18077581[28]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[28]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_a1e39e74 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[28]),
    .d(al_ccabc055[28]),
    .e(al_e45b51d9[28]),
    .o(al_c28c3a52[28]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_7d638627 (
    .a(al_e03b3126[29]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_19c0990d),
    .o(al_18077581[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_9e5fefe0 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[27]),
    .e(al_ccabc055[29]),
    .f(al_97943858[29]),
    .o(al_7b880725));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_37899172 (
    .a(al_7b880725),
    .b(al_18077581[29]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[29]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_e5add810 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[29]),
    .d(al_ccabc055[29]),
    .e(al_e45b51d9[29]),
    .o(al_c28c3a52[29]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc50fc500))
    al_64178c29 (
    .a(al_9bcd349b),
    .b(al_e03b3126[17]),
    .c(al_555b0990[0]),
    .d(al_555b0990[1]),
    .e(al_80e2c141),
    .o(al_18077581[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_c5189044 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[0]),
    .e(al_ccabc055[2]),
    .f(al_97943858[2]),
    .o(al_a34c4405));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    al_fe80e0cc (
    .a(al_a34c4405),
    .b(al_235de557),
    .c(al_4cc0b8dd),
    .d(al_1a8c7c22[2]),
    .o(al_a0c987d5));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_bd2d0dc9 (
    .a(al_a0c987d5),
    .b(al_18077581[2]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[2]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_1bee63e1 (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[2]),
    .c(al_c91705db),
    .d(al_ccabc055[2]),
    .e(al_e45b51d9[2]),
    .o(al_c28c3a52[2]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_6dc67651 (
    .a(al_e03b3126[30]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_cacb44c4),
    .o(al_18077581[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_77f1e29c (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[28]),
    .e(al_ccabc055[30]),
    .f(al_97943858[30]),
    .o(al_23658752));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_92b01270 (
    .a(al_23658752),
    .b(al_235de557),
    .c(al_9c55c5c3),
    .o(al_e9a9157c));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_d73da2b7 (
    .a(al_e9a9157c),
    .b(al_18077581[30]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[30]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_9be7e933 (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[30]),
    .c(al_c91705db),
    .d(al_ccabc055[30]),
    .e(al_e45b51d9[30]),
    .o(al_c28c3a52[30]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_4ee5968 (
    .a(al_e03b3126[31]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_14b732b9),
    .o(al_18077581[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*D)*~(E*B)*~(C*A))"),
    .INIT(64'h0013005f13135f5f))
    al_a9320bf6 (
    .a(al_ee8b2558),
    .b(al_be8ea5e1),
    .c(al_4cc0b8dd),
    .d(al_7610b7fc),
    .e(al_ccabc055[31]),
    .f(al_97943858[31]),
    .o(al_10df355f));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    al_8ec5af1b (
    .a(al_10df355f),
    .b(al_d19b9f6b),
    .c(al_35d85285[29]),
    .o(al_ed766401));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_3ba5d7d4 (
    .a(al_ed766401),
    .b(al_18077581[31]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[31]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_1cb35d3d (
    .a(al_9176d089),
    .b(al_be8ea5e1),
    .o(al_98ab69b8));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_96497a5c (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[31]),
    .c(al_c91705db),
    .d(al_ccabc055[31]),
    .e(al_e45b51d9[31]),
    .o(al_c28c3a52[31]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_5c0d1ccf (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[3]),
    .c(al_c91705db),
    .d(al_ccabc055[3]),
    .e(al_e45b51d9[3]),
    .o(al_c28c3a52[3]));
  AL_MAP_LUT4 #(
    .EQN("(A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*C*D)"),
    .INIT(16'h8380))
    al_7da1c5f4 (
    .a(al_e03b3126[19]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_5df930ee),
    .o(al_18077581[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_bd50c77c (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[2]),
    .e(al_ccabc055[4]),
    .f(al_97943858[4]),
    .o(al_7095ffb4));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_8556c2fa (
    .a(al_7095ffb4),
    .b(al_235de557),
    .o(al_e0306332));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_54ea848d (
    .a(al_e0306332),
    .b(al_18077581[4]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[4]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_2143c67a (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[4]),
    .c(al_c91705db),
    .d(al_ccabc055[4]),
    .e(al_e45b51d9[4]),
    .o(al_c28c3a52[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_1f42c5dc (
    .a(al_555b0990[0]),
    .b(al_555b0990[1]),
    .c(al_8e267e24),
    .o(al_18077581[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_4d57b23c (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[3]),
    .e(al_ccabc055[5]),
    .f(al_97943858[5]),
    .o(al_75b09ba0));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_67374afd (
    .a(al_75b09ba0),
    .b(al_18077581[5]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[5]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_8a309487 (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[5]),
    .d(al_ccabc055[5]),
    .e(al_e45b51d9[5]),
    .o(al_c28c3a52[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_c2c48a6b (
    .a(al_555b0990[0]),
    .b(al_555b0990[1]),
    .c(al_e163f204),
    .o(al_18077581[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_82656f8c (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[4]),
    .e(al_ccabc055[6]),
    .f(al_97943858[6]),
    .o(al_37698acd));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_1fac11b0 (
    .a(al_37698acd),
    .b(al_9c55c5c3),
    .o(al_bb5767ca));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_a581c77e (
    .a(al_bb5767ca),
    .b(al_18077581[6]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_9210d070 (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[6]),
    .c(al_c91705db),
    .d(al_ccabc055[6]),
    .e(al_e45b51d9[6]),
    .o(al_c28c3a52[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_50d5dfcd (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[7]),
    .c(al_c91705db),
    .d(al_ccabc055[7]),
    .e(al_e45b51d9[7]),
    .o(al_c28c3a52[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_13c8b0a7 (
    .a(al_555b0990[0]),
    .b(al_555b0990[1]),
    .c(al_a35cf148),
    .o(al_18077581[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_a4e8ae86 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[6]),
    .e(al_ccabc055[8]),
    .f(al_97943858[8]),
    .o(al_26af78f7));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_750fb4c1 (
    .a(al_26af78f7),
    .b(al_18077581[8]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)*~(A)+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*~(A)+~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*C*A+(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C*A)"),
    .INIT(32'hf5b1e4a0))
    al_4b186bea (
    .a(al_98ab69b8),
    .b(al_c91705db),
    .c(al_3bdbe1c8[8]),
    .d(al_ccabc055[8]),
    .e(al_e45b51d9[8]),
    .o(al_c28c3a52[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_a694b1cc (
    .a(al_555b0990[0]),
    .b(al_555b0990[1]),
    .c(al_728c73ac),
    .o(al_18077581[9]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_ab5a1118 (
    .a(al_d19b9f6b),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_35d85285[7]),
    .e(al_ccabc055[9]),
    .f(al_97943858[9]),
    .o(al_92fd4928));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5acf3d09 (
    .a(al_92fd4928),
    .b(al_235de557),
    .o(al_29a1a38f));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_72456112 (
    .a(al_29a1a38f),
    .b(al_18077581[9]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[9]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*~(B)*~(A)+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*~(A)+~((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C))*B*A+(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)*B*A)"),
    .INIT(32'hdd8dd888))
    al_4092f5f (
    .a(al_98ab69b8),
    .b(al_3bdbe1c8[9]),
    .c(al_c91705db),
    .d(al_ccabc055[9]),
    .e(al_e45b51d9[9]),
    .o(al_c28c3a52[9]));
  AL_DFF_X al_ebd86703 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9eda716),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da7f07ab));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e28d6f3b (
    .a(al_70d8b4ee),
    .b(al_3bdbe1c8[11]),
    .c(al_da7f07ab),
    .o(al_9eda716));
  AL_DFF_X al_292b32ac (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_29632809),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa37cfdb));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2ce18613 (
    .a(al_70d8b4ee),
    .b(al_3bdbe1c8[3]),
    .c(al_aa37cfdb),
    .o(al_29632809));
  AL_DFF_X al_6b8552a2 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e9c55e9a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_172eec6a));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_8d3bbce1 (
    .a(al_9176d089),
    .b(al_804ebeec),
    .o(al_70d8b4ee));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_21bc9e62 (
    .a(al_70d8b4ee),
    .b(al_3bdbe1c8[7]),
    .c(al_172eec6a),
    .o(al_e9c55e9a));
  AL_DFF_X al_a75be8d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_abe3d564),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8869249d));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    al_a9c08d36 (
    .a(al_9176d089),
    .b(al_3bdbe1c8[3]),
    .c(al_92eee380),
    .d(al_809b319),
    .o(al_8de27684));
  AL_DFF_X al_2e75404f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8de27684),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3697c94f));
  AL_DFF_X al_47ec0c00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_384c501e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1a600b6));
  AL_MAP_LUT4 #(
    .EQN("(A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*C*D)"),
    .INIT(16'h8380))
    al_3534d599 (
    .a(al_e03b3126[18]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_1e979a01),
    .o(al_18077581[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(D*B)*~(E*A))"),
    .INIT(64'h0105030f115533ff))
    al_9daeb86a (
    .a(al_be8ea5e1),
    .b(al_4cc0b8dd),
    .c(al_7610b7fc),
    .d(al_1a8c7c22[3]),
    .e(al_ccabc055[3]),
    .f(al_97943858[3]),
    .o(al_7b361041));
  AL_MAP_LUT6 #(
    .EQN("(~(F*E)*~(C*B)*~(D*A))"),
    .INIT(64'h0000153f153f153f))
    al_5e0887af (
    .a(al_aa37cfdb),
    .b(al_ac1a4f11),
    .c(al_e9897485),
    .d(al_804ebeec),
    .e(al_d19b9f6b),
    .f(al_35d85285[1]),
    .o(al_3d3ab166));
  AL_MAP_LUT5 #(
    .EQN("(~D*B*A*~(E*C))"),
    .INIT(32'h00080088))
    al_6ed7bb7c (
    .a(al_7b361041),
    .b(al_3d3ab166),
    .c(al_3697c94f),
    .d(al_235de557),
    .e(al_809b319),
    .o(al_1d8052bb));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_74e2642e (
    .a(al_1d8052bb),
    .b(al_18077581[3]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[3]));
  AL_MAP_LUT6 #(
    .EQN("(((E*C)*~(F)*~(D)+(E*C)*F*~(D)+~((E*C))*F*D+(E*C)*F*D)*~(B)*~(A)+((E*C)*~(F)*~(D)+(E*C)*F*~(D)+~((E*C))*F*D+(E*C)*F*D)*B*~(A)+~(((E*C)*~(F)*~(D)+(E*C)*F*~(D)+~((E*C))*F*D+(E*C)*F*D))*B*A+((E*C)*~(F)*~(D)+(E*C)*F*~(D)+~((E*C))*F*D+(E*C)*F*D)*B*A)"),
    .INIT(64'hddd8dd8888d88888))
    al_80f8cd99 (
    .a(al_4989df73),
    .b(al_3bdbe1c8[3]),
    .c(al_c91705db),
    .d(al_53cc722d),
    .e(al_ac1a4f11),
    .f(al_4d792cee),
    .o(al_74d8fce0));
  AL_DFF_X al_83e2843e (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_74d8fce0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1a4f11));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_3ca437a9 (
    .a(al_555b0990[0]),
    .b(al_555b0990[1]),
    .c(al_a6e0ed04),
    .o(al_18077581[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*D)*~(C*B)*~(E*A))"),
    .INIT(64'h0015003f15153f3f))
    al_9edddd3f (
    .a(al_a1a600b6),
    .b(al_4d792cee),
    .c(al_e9897485),
    .d(al_be8ea5e1),
    .e(al_809b319),
    .f(al_ccabc055[7]),
    .o(al_1b41bac1));
  AL_MAP_LUT6 #(
    .EQN("(~(F*D)*~(E*C)*~(B*A))"),
    .INIT(64'h0007007707077777))
    al_29f4f5a3 (
    .a(al_172eec6a),
    .b(al_804ebeec),
    .c(al_d19b9f6b),
    .d(al_7610b7fc),
    .e(al_35d85285[5]),
    .f(al_97943858[7]),
    .o(al_7242df1f));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_8039f326 (
    .a(al_1b41bac1),
    .b(al_7242df1f),
    .c(al_235de557),
    .o(al_83268b9b));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_2acc275a (
    .a(al_83268b9b),
    .b(al_18077581[7]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(~D*~(E*~(F)*~(C)+E*F*~(C)+~(E)*F*C+E*F*C))*~(B)*~(A)+~(~D*~(E*~(F)*~(C)+E*F*~(C)+~(E)*F*C+E*F*C))*B*~(A)+~(~(~D*~(E*~(F)*~(C)+E*F*~(C)+~(E)*F*C+E*F*C)))*B*A+~(~D*~(E*~(F)*~(C)+E*F*~(C)+~(E)*F*C+E*F*C))*B*A)"),
    .INIT(64'hddddddd8dd8ddd88))
    al_8c47276 (
    .a(al_4989df73),
    .b(al_3bdbe1c8[7]),
    .c(al_c91705db),
    .d(al_53cc722d),
    .e(al_ac1a4f11),
    .f(al_4d792cee),
    .o(al_c1679159));
  AL_DFF_X al_32b211c3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1679159),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4d792cee));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_9227596 (
    .a(al_555b0990[0]),
    .b(al_555b0990[1]),
    .c(al_fdf9f0dc),
    .o(al_18077581[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(D*B)*~(E*A))"),
    .INIT(64'h0105030f115533ff))
    al_832eebbf (
    .a(al_e9897485),
    .b(al_d19b9f6b),
    .c(al_7610b7fc),
    .d(al_35d85285[9]),
    .e(al_12792818[0]),
    .f(al_97943858[11]),
    .o(al_48dfd35c));
  AL_MAP_LUT6 #(
    .EQN("(~(F*D)*~(E*B)*~(C*A))"),
    .INIT(64'h0013005f13135f5f))
    al_c25521a4 (
    .a(al_da7f07ab),
    .b(al_8869249d),
    .c(al_804ebeec),
    .d(al_be8ea5e1),
    .e(al_809b319),
    .f(al_ccabc055[11]),
    .o(al_1de941c8));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_c3259199 (
    .a(al_48dfd35c),
    .b(al_1de941c8),
    .c(al_235de557),
    .o(al_5f34afe1));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_1498ccbb (
    .a(al_5f34afe1),
    .b(al_18077581[11]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[11]));
  AL_MAP_LUT5 #(
    .EQN("((~D*~(~E*C))*~(B)*~(A)+(~D*~(~E*C))*B*~(A)+~((~D*~(~E*C)))*B*A+(~D*~(~E*C))*B*A)"),
    .INIT(32'h88dd888d))
    al_f0105bd (
    .a(al_4989df73),
    .b(al_3bdbe1c8[11]),
    .c(al_c91705db),
    .d(al_53cc722d),
    .e(al_12792818[0]),
    .o(al_591b5570[0]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_e6049636 (
    .a(al_bb6625de[1]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_b5bf2603),
    .o(al_18077581[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(D*B)*~(E*A))"),
    .INIT(64'h0105030f115533ff))
    al_45f0c3fe (
    .a(al_e9897485),
    .b(al_be8ea5e1),
    .c(al_7610b7fc),
    .d(al_ccabc055[12]),
    .e(al_12792818[1]),
    .f(al_97943858[12]),
    .o(al_fdd40d67));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    al_9d29739b (
    .a(al_fdd40d67),
    .b(al_235de557),
    .c(al_d19b9f6b),
    .d(al_35d85285[10]),
    .o(al_63c14fc));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1dcc))
    al_79e9d6b5 (
    .a(al_63c14fc),
    .b(al_18077581[12]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_3bdbe1c8[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_73170fb0 (
    .a(al_5a744f0f),
    .b(al_b211b12d),
    .c(al_39cb3b56),
    .o(al_9176d089));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_8c9ef44b (
    .a(al_9176d089),
    .b(al_e9897485),
    .o(al_4989df73));
  AL_MAP_LUT5 #(
    .EQN("((~D*~(~E*C))*~(B)*~(A)+(~D*~(~E*C))*B*~(A)+~((~D*~(~E*C)))*B*A+(~D*~(~E*C))*B*A)"),
    .INIT(32'h88dd888d))
    al_f0945b02 (
    .a(al_4989df73),
    .b(al_3bdbe1c8[12]),
    .c(al_c91705db),
    .d(al_53cc722d),
    .e(al_12792818[1]),
    .o(al_591b5570[1]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*~B))"),
    .INIT(16'ha080))
    al_fdb68f89 (
    .a(al_3f1d46e5),
    .b(al_5a744f0f),
    .c(al_c197c567),
    .d(al_16745a5f),
    .o(al_a63110e1));
  AL_DFF_X al_9b5f8bd4 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a63110e1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16745a5f));
  AL_MAP_LUT5 #(
    .EQN("(C*A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))"),
    .INIT(32'ha0208000))
    al_a152b297 (
    .a(al_3f1d46e5),
    .b(al_bb0cd305),
    .c(al_c197c567),
    .d(al_16745a5f),
    .e(al_f5b6a552),
    .o(al_75e66ec7));
  AL_DFF_X al_f93c5848 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_75e66ec7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5b6a552));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_37fe08c1 (
    .a(al_3f1d46e5),
    .b(al_c197c567),
    .c(al_f5b6a552),
    .o(al_d119a42b));
  AL_DFF_X al_84d03779 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d119a42b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2a43721c));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_e6a740c (
    .a(al_6fd79ca[0]),
    .b(al_e4d248a4),
    .c(al_43722bf9[0]),
    .d(al_9bf95cff[0]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_a6d94861 (
    .a(al_6fd79ca[10]),
    .b(al_e4d248a4),
    .c(al_43722bf9[10]),
    .d(al_9bf95cff[10]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[10]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_e91cd7f1 (
    .a(al_6fd79ca[11]),
    .b(al_e4d248a4),
    .c(al_43722bf9[11]),
    .d(al_9bf95cff[11]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[11]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_7ce0d1e3 (
    .a(al_6fd79ca[12]),
    .b(al_e4d248a4),
    .c(al_43722bf9[12]),
    .d(al_9bf95cff[12]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[12]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_12093b7d (
    .a(al_6fd79ca[13]),
    .b(al_e4d248a4),
    .c(al_43722bf9[13]),
    .d(al_9bf95cff[13]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[13]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_9b244e62 (
    .a(al_6fd79ca[14]),
    .b(al_e4d248a4),
    .c(al_43722bf9[14]),
    .d(al_9bf95cff[14]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[14]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_befee68a (
    .a(al_6fd79ca[15]),
    .b(al_e4d248a4),
    .c(al_43722bf9[15]),
    .d(al_9bf95cff[15]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[15]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_7981d068 (
    .a(al_6fd79ca[16]),
    .b(al_e4d248a4),
    .c(al_43722bf9[16]),
    .d(al_9bf95cff[16]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[16]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_14c9247d (
    .a(al_6fd79ca[17]),
    .b(al_e4d248a4),
    .c(al_43722bf9[17]),
    .d(al_9bf95cff[17]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[17]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_43edc248 (
    .a(al_6fd79ca[18]),
    .b(al_e4d248a4),
    .c(al_43722bf9[18]),
    .d(al_9bf95cff[18]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[18]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_51115421 (
    .a(al_6fd79ca[19]),
    .b(al_e4d248a4),
    .c(al_43722bf9[19]),
    .d(al_9bf95cff[19]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[19]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_d0cbb5be (
    .a(al_6fd79ca[1]),
    .b(al_e4d248a4),
    .c(al_43722bf9[1]),
    .d(al_9bf95cff[1]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_f8d5d505 (
    .a(al_6fd79ca[20]),
    .b(al_e4d248a4),
    .c(al_43722bf9[20]),
    .d(al_9bf95cff[20]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[20]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_f4782a8c (
    .a(al_6fd79ca[21]),
    .b(al_e4d248a4),
    .c(al_43722bf9[21]),
    .d(al_9bf95cff[21]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[21]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_e5945804 (
    .a(al_6fd79ca[22]),
    .b(al_e4d248a4),
    .c(al_43722bf9[22]),
    .d(al_9bf95cff[22]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[22]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_6d3ae833 (
    .a(al_6fd79ca[23]),
    .b(al_e4d248a4),
    .c(al_43722bf9[23]),
    .d(al_9bf95cff[23]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[23]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_4969a841 (
    .a(al_6fd79ca[24]),
    .b(al_e4d248a4),
    .c(al_43722bf9[24]),
    .d(al_9bf95cff[24]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[24]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_e2fd5d13 (
    .a(al_6fd79ca[25]),
    .b(al_e4d248a4),
    .c(al_43722bf9[25]),
    .d(al_9bf95cff[25]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[25]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_3411cc4c (
    .a(al_6fd79ca[26]),
    .b(al_e4d248a4),
    .c(al_43722bf9[26]),
    .d(al_9bf95cff[26]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[26]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_2cc31029 (
    .a(al_6fd79ca[27]),
    .b(al_e4d248a4),
    .c(al_43722bf9[27]),
    .d(al_9bf95cff[27]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[27]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_2ff5e34a (
    .a(al_6fd79ca[28]),
    .b(al_e4d248a4),
    .c(al_43722bf9[28]),
    .d(al_9bf95cff[28]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[28]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_7f21736b (
    .a(al_6fd79ca[29]),
    .b(al_e4d248a4),
    .c(al_43722bf9[29]),
    .d(al_9bf95cff[29]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[29]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_a1184e83 (
    .a(al_6fd79ca[2]),
    .b(al_e4d248a4),
    .c(al_43722bf9[2]),
    .d(al_9bf95cff[2]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[2]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_e79d8a4c (
    .a(al_6fd79ca[30]),
    .b(al_e4d248a4),
    .c(al_43722bf9[30]),
    .d(al_9bf95cff[30]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[30]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_68098ee8 (
    .a(al_6fd79ca[31]),
    .b(al_e4d248a4),
    .c(al_43722bf9[31]),
    .d(al_9bf95cff[31]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[31]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_93b1018b (
    .a(al_6fd79ca[3]),
    .b(al_e4d248a4),
    .c(al_43722bf9[3]),
    .d(al_9bf95cff[3]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_d7f33f0d (
    .a(al_6fd79ca[4]),
    .b(al_e4d248a4),
    .c(al_43722bf9[4]),
    .d(al_9bf95cff[4]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[4]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_47947ae6 (
    .a(al_6fd79ca[5]),
    .b(al_e4d248a4),
    .c(al_43722bf9[5]),
    .d(al_9bf95cff[5]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[5]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_dfef7ee7 (
    .a(al_6fd79ca[6]),
    .b(al_e4d248a4),
    .c(al_43722bf9[6]),
    .d(al_9bf95cff[6]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[6]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_a4fb4ad0 (
    .a(al_6fd79ca[7]),
    .b(al_e4d248a4),
    .c(al_43722bf9[7]),
    .d(al_9bf95cff[7]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[7]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_da4b8c03 (
    .a(al_6fd79ca[8]),
    .b(al_e4d248a4),
    .c(al_43722bf9[8]),
    .d(al_9bf95cff[8]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[8]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*~(D)*~(B)+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*~(B)+~((C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E))*D*B+(C*~(A)*~(E)+C*A*~(E)+~(C)*A*E+C*A*E)*D*B)"),
    .INIT(32'hee22fc30))
    al_c35d6b45 (
    .a(al_6fd79ca[9]),
    .b(al_e4d248a4),
    .c(al_43722bf9[9]),
    .d(al_9bf95cff[9]),
    .e(al_c0a7a5f),
    .o(al_d610ac57[9]));
  AL_DFF_X al_131b31b0 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c3006fde),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afb86315));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_adb5302d (
    .a(al_4cb17b0d),
    .b(al_afb86315),
    .o(al_c3006fde));
  AL_DFF_X al_e05d7720 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f325673f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_67635cb3));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*B*C*D)"),
    .INIT(16'h44ec))
    al_f2fc53d5 (
    .a(al_2c4c1ef7),
    .b(al_67635cb3),
    .c(al_25fbce42[50]),
    .d(al_25fbce42[58]),
    .o(al_f325673f));
  AL_MAP_LUT5 #(
    .EQN("(~(~(~D*C)*~B)*~(E*A))"),
    .INIT(32'h4454ccfc))
    al_45a3beb1 (
    .a(al_2c4c1ef7),
    .b(al_8c0460e8),
    .c(al_6893b11d),
    .d(al_52c6af0a),
    .e(al_25fbce42[57]),
    .o(al_76e89bee));
  AL_DFF_X al_798d9b06 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_76e89bee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c0460e8));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_806f5351 (
    .a(al_a27f756f),
    .b(al_25fbce42[2]),
    .o(al_2c4c1ef7));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(C*~B*~(~E*~D)))"),
    .INIT(32'h45454555))
    al_8da401b8 (
    .a(al_e379ebb5),
    .b(al_f6cd735f),
    .c(al_69807e37),
    .d(al_f49992c3),
    .e(al_c73c0ba3),
    .o(al_2482626f));
  AL_MAP_LUT5 #(
    .EQN("~(B*(~(A)*~(C)*~(D)*~(E)+A*~(C)*~(D)*~(E)+~(A)*~(C)*D*~(E)+~(A)*~(C)*~(D)*E+A*~(C)*~(D)*E+A*C*~(D)*E+~(A)*~(C)*D*E+A*~(C)*D*E+A*C*D*E))"),
    .INIT(32'h7373fbf3))
    al_ea2e7111 (
    .a(al_2c4c1ef7),
    .b(al_2482626f),
    .c(al_6893b11d),
    .d(al_25fbce42[49]),
    .e(al_25fbce42[57]),
    .o(al_30c029d2));
  AL_DFF_X al_922bf2c1 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_30c029d2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6893b11d));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(C*~(D*A)))"),
    .INIT(16'hdcfc))
    al_c883695a (
    .a(al_2c4c1ef7),
    .b(al_e379ebb5),
    .c(al_6f63d541),
    .d(al_25fbce42[57]),
    .o(al_8805aafa));
  AL_DFF_X al_684674bf (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8805aafa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f63d541));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~D*~C*~B*A)"),
    .INIT(32'hfffffffd))
    al_c633aea3 (
    .a(al_f6cd735f),
    .b(al_f49992c3),
    .c(al_523cde28),
    .d(al_501dbbdf),
    .e(al_c0a7a5f),
    .o(al_8f2c85dc));
  AL_DFF_X al_f1605192 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8f2c85dc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_52c6af0a));
  AL_DFF_X al_b80d6c58 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3d3aa49b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b799bc04));
  AL_DFF_X al_7ae19d02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b799bc04),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50debbc6));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*B*C*D)"),
    .INIT(16'h44ec))
    al_88886844 (
    .a(al_2c4c1ef7),
    .b(al_b799bc04),
    .c(al_25fbce42[48]),
    .d(al_25fbce42[56]),
    .o(al_3d3aa49b));
  AL_DFF_X al_8a7de15d (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8e7f80da),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_69807e37));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c9e18ae8 (
    .a(al_2c4c1ef7),
    .b(al_69807e37),
    .c(al_25fbce42[36]),
    .o(al_8e7f80da));
  AL_DFF_X al_182451a0 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_5493f072),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b3a31b1c));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_6d789db0 (
    .a(al_4ed450cb),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[10]),
    .e(al_683f5875[8]),
    .o(al_40185430[10]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_ca10fa69 (
    .a(al_667db93d),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[11]),
    .e(al_683f5875[9]),
    .o(al_40185430[11]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_2f099f0c (
    .a(al_fb26226a),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[12]),
    .e(al_683f5875[10]),
    .o(al_40185430[12]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_ce560b87 (
    .a(al_c4d4b7f5),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[13]),
    .e(al_683f5875[11]),
    .o(al_40185430[13]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_cad40b49 (
    .a(al_13708b94),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[14]),
    .e(al_683f5875[12]),
    .o(al_40185430[14]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_849a86de (
    .a(al_8cb8f5f5),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[15]),
    .e(al_683f5875[13]),
    .o(al_40185430[15]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_32809a07 (
    .a(al_c5cc2f9b),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[16]),
    .e(al_683f5875[14]),
    .o(al_40185430[16]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_df02e6fb (
    .a(al_c048f5a0),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[17]),
    .e(al_683f5875[15]),
    .o(al_40185430[17]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_fb4aa692 (
    .a(al_c6cd8be8),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[18]),
    .e(al_683f5875[16]),
    .o(al_40185430[18]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_a5d6f42b (
    .a(al_31822056),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[19]),
    .e(al_683f5875[17]),
    .o(al_40185430[19]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_a05d01df (
    .a(al_6e8dae0d),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[20]),
    .e(al_683f5875[18]),
    .o(al_40185430[20]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_a01b6ba7 (
    .a(al_f76f8d54),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[21]),
    .e(al_683f5875[19]),
    .o(al_40185430[21]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_421a1daa (
    .a(al_825438f5),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[22]),
    .e(al_683f5875[20]),
    .o(al_40185430[22]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_ee60c34 (
    .a(al_ab46d2b9),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[23]),
    .e(al_683f5875[21]),
    .o(al_40185430[23]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_9d5308a1 (
    .a(al_d33dd538),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[24]),
    .e(al_683f5875[22]),
    .o(al_40185430[24]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_2e65cc88 (
    .a(al_b62de081),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[25]),
    .e(al_683f5875[23]),
    .o(al_40185430[25]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_7dee996f (
    .a(al_447f0158),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[26]),
    .e(al_683f5875[24]),
    .o(al_40185430[26]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_307c033e (
    .a(al_a0670bff),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[27]),
    .e(al_683f5875[25]),
    .o(al_40185430[27]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_6bfa1c58 (
    .a(al_74973e72),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[28]),
    .e(al_683f5875[26]),
    .o(al_40185430[28]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_2310e8b7 (
    .a(al_cae3c642),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[29]),
    .e(al_683f5875[27]),
    .o(al_40185430[29]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_d80b7568 (
    .a(al_3db1ed2d),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[2]),
    .e(al_683f5875[0]),
    .o(al_40185430[2]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_85f3e9fa (
    .a(al_ac5b8836),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[30]),
    .e(al_683f5875[28]),
    .o(al_40185430[30]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_7a69e98b (
    .a(al_9bb19ed8),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[31]),
    .e(al_683f5875[29]),
    .o(al_40185430[31]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_3eb9e1b (
    .a(al_e9dadc09),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[3]),
    .e(al_683f5875[1]),
    .o(al_40185430[3]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_ad129a01 (
    .a(al_3be09bce),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[4]),
    .e(al_683f5875[2]),
    .o(al_40185430[4]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_6467d953 (
    .a(al_8773b31),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[5]),
    .e(al_683f5875[3]),
    .o(al_40185430[5]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_fd9e1266 (
    .a(al_640ea1c6),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[6]),
    .e(al_683f5875[4]),
    .o(al_40185430[6]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_d7da2325 (
    .a(al_4e819ed5),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[7]),
    .e(al_683f5875[5]),
    .o(al_40185430[7]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_f7a1a26b (
    .a(al_2418b5af),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[8]),
    .e(al_683f5875[6]),
    .o(al_40185430[8]));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*~(D)*~(C)+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*~(C)+~((~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B))*D*C+(~A*~(E)*~(B)+~A*E*~(B)+~(~A)*E*B+~A*E*B)*D*C)"),
    .INIT(32'hfd0df101))
    al_114f0464 (
    .a(al_4a696460),
    .b(al_fa66b6a3),
    .c(al_48d2ef94),
    .d(al_8c9327d6[9]),
    .e(al_683f5875[7]),
    .o(al_40185430[9]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(~C*B*A))"),
    .INIT(16'hff08))
    al_301baac2 (
    .a(al_a25a6119),
    .b(al_c83b3308),
    .c(al_66ffb9),
    .d(al_48d2ef94),
    .o(al_6897cc6d));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~(~C*B*A)))"),
    .INIT(32'h00ff0008))
    al_7abcec59 (
    .a(al_a25a6119),
    .b(al_c83b3308),
    .c(al_66ffb9),
    .d(iBusAhb_HREADY),
    .e(al_48d2ef94),
    .o(al_7408b2ea));
  AL_DFF_X al_7c1170f5 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_7408b2ea),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48d2ef94));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_8b05203 (
    .a(al_48d2ef94),
    .o(al_766b3b75));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_9f2e07c3 (
    .a(1'b0),
    .o({al_10ccc4a2,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c6771808 (
    .a(al_a16ef20a[1]),
    .b(al_24a3e858),
    .c(al_10ccc4a2),
    .o({al_7fea1a88,al_b24d99c7[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7844c7cc (
    .a(al_a16ef20a[2]),
    .b(al_6515336d[2]),
    .c(al_7fea1a88),
    .o({al_90ed329,al_b24d99c7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ff5f2dcb (
    .a(al_a16ef20a[3]),
    .b(1'b0),
    .c(al_90ed329),
    .o({al_6d5a6293,al_b24d99c7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_72840809 (
    .a(al_a16ef20a[4]),
    .b(1'b0),
    .c(al_6d5a6293),
    .o({al_aa88d0b2,al_b24d99c7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e70bb85a (
    .a(al_a16ef20a[5]),
    .b(1'b0),
    .c(al_aa88d0b2),
    .o({al_6ecad7e7,al_b24d99c7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c0755da (
    .a(al_a16ef20a[6]),
    .b(1'b0),
    .c(al_6ecad7e7),
    .o({al_42d0475,al_b24d99c7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4fe7e2af (
    .a(al_a16ef20a[7]),
    .b(1'b0),
    .c(al_42d0475),
    .o({al_927566f,al_b24d99c7[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9a6823a2 (
    .a(al_a16ef20a[8]),
    .b(1'b0),
    .c(al_927566f),
    .o({al_18e9bd9b,al_b24d99c7[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b4911995 (
    .a(al_a16ef20a[9]),
    .b(1'b0),
    .c(al_18e9bd9b),
    .o({al_e2f2e915,al_b24d99c7[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bcc5ba40 (
    .a(al_a16ef20a[10]),
    .b(1'b0),
    .c(al_e2f2e915),
    .o({al_d0a81721,al_b24d99c7[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7e89c44e (
    .a(al_a16ef20a[11]),
    .b(1'b0),
    .c(al_d0a81721),
    .o({al_f529ac86,al_b24d99c7[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f87055a5 (
    .a(al_a16ef20a[12]),
    .b(1'b0),
    .c(al_f529ac86),
    .o({al_13bd3caf,al_b24d99c7[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b3bbc1c1 (
    .a(al_a16ef20a[13]),
    .b(1'b0),
    .c(al_13bd3caf),
    .o({al_52ea8e26,al_b24d99c7[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_89fcdf09 (
    .a(al_a16ef20a[14]),
    .b(1'b0),
    .c(al_52ea8e26),
    .o({al_f0a4b18b,al_b24d99c7[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cdf43596 (
    .a(al_a16ef20a[15]),
    .b(1'b0),
    .c(al_f0a4b18b),
    .o({al_1e389db1,al_b24d99c7[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d91f0f24 (
    .a(al_a16ef20a[16]),
    .b(1'b0),
    .c(al_1e389db1),
    .o({al_123d8e5f,al_b24d99c7[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5e9eab80 (
    .a(al_a16ef20a[17]),
    .b(1'b0),
    .c(al_123d8e5f),
    .o({al_a241616a,al_b24d99c7[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bd6fb13b (
    .a(al_a16ef20a[18]),
    .b(1'b0),
    .c(al_a241616a),
    .o({al_8e70d65a,al_b24d99c7[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_238009de (
    .a(al_a16ef20a[19]),
    .b(1'b0),
    .c(al_8e70d65a),
    .o({al_45ceabc3,al_b24d99c7[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a6084fa6 (
    .a(al_a16ef20a[20]),
    .b(1'b0),
    .c(al_45ceabc3),
    .o({al_19e34f5d,al_b24d99c7[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6bffe9df (
    .a(al_a16ef20a[21]),
    .b(1'b0),
    .c(al_19e34f5d),
    .o({al_9a97f855,al_b24d99c7[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7dec2c74 (
    .a(al_a16ef20a[22]),
    .b(1'b0),
    .c(al_9a97f855),
    .o({al_edcbe33d,al_b24d99c7[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_95457dcb (
    .a(al_a16ef20a[23]),
    .b(1'b0),
    .c(al_edcbe33d),
    .o({al_91a72f10,al_b24d99c7[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cf321750 (
    .a(al_a16ef20a[24]),
    .b(1'b0),
    .c(al_91a72f10),
    .o({al_a59daeb4,al_b24d99c7[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d116c1e1 (
    .a(al_a16ef20a[25]),
    .b(1'b0),
    .c(al_a59daeb4),
    .o({al_781bb51f,al_b24d99c7[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d584ec61 (
    .a(al_a16ef20a[26]),
    .b(1'b0),
    .c(al_781bb51f),
    .o({al_d4ff0ad3,al_b24d99c7[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_10cc5bef (
    .a(al_a16ef20a[27]),
    .b(1'b0),
    .c(al_d4ff0ad3),
    .o({al_ffb1962,al_b24d99c7[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dd304edd (
    .a(al_a16ef20a[28]),
    .b(1'b0),
    .c(al_ffb1962),
    .o({al_443f5c3a,al_b24d99c7[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ecfc1826 (
    .a(al_a16ef20a[29]),
    .b(1'b0),
    .c(al_443f5c3a),
    .o({al_d2147867,al_b24d99c7[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dba67d93 (
    .a(al_a16ef20a[30]),
    .b(1'b0),
    .c(al_d2147867),
    .o({al_1e7955bd,al_b24d99c7[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_54184c3b (
    .a(al_a16ef20a[31]),
    .b(1'b0),
    .c(al_1e7955bd),
    .o({open_n7,al_b24d99c7[30]}));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_dd4ab82c (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[8]),
    .d(al_46ea2d9f[10]),
    .e(al_ccabc055[10]),
    .f(al_2cd19c12),
    .o(al_4ed450cb));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_927c1450 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_4ed450cb),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[10]),
    .f(al_b24d99c7[9]),
    .o(al_bde0dc95[10]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_89551897 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[9]),
    .d(al_46ea2d9f[11]),
    .e(al_ccabc055[11]),
    .f(al_cc989ac9),
    .o(al_667db93d));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_76b3a3c9 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_667db93d),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[11]),
    .f(al_b24d99c7[10]),
    .o(al_bde0dc95[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_fa079c51 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[10]),
    .d(al_46ea2d9f[12]),
    .e(al_ccabc055[12]),
    .f(al_1953385a),
    .o(al_fb26226a));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_4cb70082 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_fb26226a),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[12]),
    .f(al_b24d99c7[11]),
    .o(al_bde0dc95[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_19e59acc (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[11]),
    .d(al_46ea2d9f[13]),
    .e(al_ccabc055[13]),
    .f(al_be6e0599),
    .o(al_c4d4b7f5));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_19cab682 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_c4d4b7f5),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[13]),
    .f(al_b24d99c7[12]),
    .o(al_bde0dc95[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_1c459f26 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[12]),
    .d(al_46ea2d9f[14]),
    .e(al_ccabc055[14]),
    .f(al_afe5948f),
    .o(al_13708b94));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_683b858b (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_13708b94),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[14]),
    .f(al_b24d99c7[13]),
    .o(al_bde0dc95[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_4bf40637 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[13]),
    .d(al_46ea2d9f[15]),
    .e(al_ccabc055[15]),
    .f(al_d1fc8906),
    .o(al_8cb8f5f5));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_c2a407a5 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_8cb8f5f5),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[15]),
    .f(al_b24d99c7[14]),
    .o(al_bde0dc95[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_22a617e4 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[14]),
    .d(al_46ea2d9f[16]),
    .e(al_ccabc055[16]),
    .f(al_9df5b848),
    .o(al_c5cc2f9b));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_67fb52af (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_c5cc2f9b),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[16]),
    .f(al_b24d99c7[15]),
    .o(al_bde0dc95[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_e6167345 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[15]),
    .d(al_46ea2d9f[17]),
    .e(al_ccabc055[17]),
    .f(al_afd990ff),
    .o(al_c048f5a0));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_696f62a5 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_c048f5a0),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[17]),
    .f(al_b24d99c7[16]),
    .o(al_bde0dc95[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_d8f680f6 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[16]),
    .d(al_46ea2d9f[18]),
    .e(al_ccabc055[18]),
    .f(al_7bf844c2),
    .o(al_c6cd8be8));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_99814688 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_c6cd8be8),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[18]),
    .f(al_b24d99c7[17]),
    .o(al_bde0dc95[18]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_741d0df1 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[17]),
    .d(al_46ea2d9f[19]),
    .e(al_ccabc055[19]),
    .f(al_b6803a27),
    .o(al_31822056));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_fe454233 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_31822056),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[19]),
    .f(al_b24d99c7[18]),
    .o(al_bde0dc95[19]));
  AL_MAP_LUT6 #(
    .EQN("(~(E*C)*~(D*B)*~(F*A))"),
    .INIT(64'h01051155030f33ff))
    al_ee58fcf4 (
    .a(al_ee66e790),
    .b(al_1c02d8ab),
    .c(al_53cc722d),
    .d(al_46ea2d9f[1]),
    .e(al_ccabc055[1]),
    .f(al_6ae2a07d),
    .o(al_81e43d4));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((C*B))+E*F*~((C*B))+~(E)*F*(C*B)+E*F*(C*B))*~(D)*~(A)+~(E*~(F)*~((C*B))+E*F*~((C*B))+~(E)*F*(C*B)+E*F*(C*B))*D*~(A)+~(~(E*~(F)*~((C*B))+E*F*~((C*B))+~(E)*F*(C*B)+E*F*(C*B)))*D*A+~(E*~(F)*~((C*B))+E*F*~((C*B))+~(E)*F*(C*B)+E*F*(C*B))*D*A)"),
    .INIT(64'h55ff40ea15bf00aa))
    al_2fe838c3 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_3f1d46e5),
    .d(al_81e43d4),
    .e(al_a16ef20a[1]),
    .f(al_b24d99c7[0]),
    .o(al_bde0dc95[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_861e0171 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[18]),
    .d(al_46ea2d9f[20]),
    .e(al_ccabc055[20]),
    .f(al_20b06ef3),
    .o(al_6e8dae0d));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_112d0465 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_6e8dae0d),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[20]),
    .f(al_b24d99c7[19]),
    .o(al_bde0dc95[20]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_2e691b82 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[19]),
    .d(al_46ea2d9f[21]),
    .e(al_ccabc055[21]),
    .f(al_b40171bd),
    .o(al_f76f8d54));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_ee9e213 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_f76f8d54),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[21]),
    .f(al_b24d99c7[20]),
    .o(al_bde0dc95[21]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_eb4b7d92 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[20]),
    .d(al_46ea2d9f[22]),
    .e(al_ccabc055[22]),
    .f(al_42b103ed),
    .o(al_825438f5));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_ea13455 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_825438f5),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[22]),
    .f(al_b24d99c7[21]),
    .o(al_bde0dc95[22]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_2741670c (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[21]),
    .d(al_46ea2d9f[23]),
    .e(al_ccabc055[23]),
    .f(al_5a93aea7),
    .o(al_ab46d2b9));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_6321841c (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_ab46d2b9),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[23]),
    .f(al_b24d99c7[22]),
    .o(al_bde0dc95[23]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_1972a4ed (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[22]),
    .d(al_46ea2d9f[24]),
    .e(al_ccabc055[24]),
    .f(al_40d63aa3),
    .o(al_d33dd538));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_5ad118bb (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_d33dd538),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[24]),
    .f(al_b24d99c7[23]),
    .o(al_bde0dc95[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_6584cc18 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[23]),
    .d(al_46ea2d9f[25]),
    .e(al_ccabc055[25]),
    .f(al_89782fa0),
    .o(al_b62de081));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_fab9a7d0 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_b62de081),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[25]),
    .f(al_b24d99c7[24]),
    .o(al_bde0dc95[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_37455995 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[24]),
    .d(al_46ea2d9f[26]),
    .e(al_ccabc055[26]),
    .f(al_faaecf2),
    .o(al_447f0158));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_df7a9ef9 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_447f0158),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[26]),
    .f(al_b24d99c7[25]),
    .o(al_bde0dc95[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_b50f3757 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[25]),
    .d(al_46ea2d9f[27]),
    .e(al_ccabc055[27]),
    .f(al_ad2a00e5),
    .o(al_a0670bff));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_25055db1 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_a0670bff),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[27]),
    .f(al_b24d99c7[26]),
    .o(al_bde0dc95[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_19df2b0b (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[26]),
    .d(al_46ea2d9f[28]),
    .e(al_ccabc055[28]),
    .f(al_193c583f),
    .o(al_74973e72));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_65fb4c52 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_74973e72),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[28]),
    .f(al_b24d99c7[27]),
    .o(al_bde0dc95[28]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_db642f05 (
    .a(al_c795a432),
    .b(al_a8151162),
    .o(al_3f1d46e5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_be149ba1 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[27]),
    .d(al_46ea2d9f[29]),
    .e(al_ccabc055[29]),
    .f(al_a155e0b3),
    .o(al_cae3c642));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*B*~A))"),
    .INIT(16'h0b0f))
    al_9919f367 (
    .a(al_a7b01c14[2]),
    .b(al_c795a432),
    .c(al_fa66b6a3),
    .d(al_a8151162),
    .o(al_6f809586));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_5b906373 (
    .a(al_a7b01c14[2]),
    .b(al_f6cd735f),
    .c(al_8905c135),
    .o(al_e87ca79));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_3476bd36 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_cae3c642),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[29]),
    .f(al_b24d99c7[28]),
    .o(al_bde0dc95[29]));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*A*~(E*D))"),
    .INIT(32'h00080808))
    al_2ac331f0 (
    .a(al_c91705db),
    .b(al_2c3e73df),
    .c(al_ea2eaeb1),
    .d(al_cd3d5e6f),
    .e(al_501dbbdf),
    .o(al_ee66e790));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    al_585fb978 (
    .a(al_c91705db),
    .b(al_ea2eaeb1),
    .c(al_cd3d5e6f),
    .d(al_501dbbdf),
    .o(al_1c02d8ab));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_3e8ad643 (
    .a(al_ee66e790),
    .b(al_1c02d8ab),
    .o(al_8db3355a));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_408981b4 (
    .a(al_ea2eaeb1),
    .b(al_36a894af[28]),
    .c(al_36a894af[29]),
    .o(al_53cc722d));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_61a110cd (
    .a(al_ee66e790),
    .b(al_53cc722d),
    .o(al_dd37dc5d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_d614c39a (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[0]),
    .d(al_46ea2d9f[2]),
    .e(al_ccabc055[2]),
    .f(al_cc5bfca5),
    .o(al_3db1ed2d));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_e98f9861 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_3db1ed2d),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[2]),
    .f(al_b24d99c7[1]),
    .o(al_bde0dc95[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_91383909 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[28]),
    .d(al_46ea2d9f[30]),
    .e(al_ccabc055[30]),
    .f(al_89bb053a),
    .o(al_ac5b8836));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_fffaf3fd (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_ac5b8836),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[30]),
    .f(al_b24d99c7[29]),
    .o(al_bde0dc95[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_6154e029 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[29]),
    .d(al_46ea2d9f[31]),
    .e(al_ccabc055[31]),
    .f(al_4efe0c98),
    .o(al_9bb19ed8));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_945b35e5 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_9bb19ed8),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[31]),
    .f(al_b24d99c7[30]),
    .o(al_bde0dc95[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_2bc63082 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[1]),
    .d(al_46ea2d9f[3]),
    .e(al_ccabc055[3]),
    .f(al_5bcd7a0),
    .o(al_e9dadc09));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_2d7a413 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_e9dadc09),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[3]),
    .f(al_b24d99c7[2]),
    .o(al_bde0dc95[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_f22356fb (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[2]),
    .d(al_46ea2d9f[4]),
    .e(al_ccabc055[4]),
    .f(al_3ab03292),
    .o(al_3be09bce));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_210fc804 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_3be09bce),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[4]),
    .f(al_b24d99c7[3]),
    .o(al_bde0dc95[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_ac17a40c (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[3]),
    .d(al_46ea2d9f[5]),
    .e(al_ccabc055[5]),
    .f(al_22da7862),
    .o(al_8773b31));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_5eee431e (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_8773b31),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[5]),
    .f(al_b24d99c7[4]),
    .o(al_bde0dc95[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_9e7af142 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[4]),
    .d(al_46ea2d9f[6]),
    .e(al_ccabc055[6]),
    .f(al_45322fba),
    .o(al_640ea1c6));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_5f23eb55 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_640ea1c6),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[6]),
    .f(al_b24d99c7[5]),
    .o(al_bde0dc95[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_505a95cd (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[5]),
    .d(al_46ea2d9f[7]),
    .e(al_ccabc055[7]),
    .f(al_c585508d),
    .o(al_4e819ed5));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_f19864d5 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_4e819ed5),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[7]),
    .f(al_b24d99c7[6]),
    .o(al_bde0dc95[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_c2bf6cc5 (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[6]),
    .d(al_46ea2d9f[8]),
    .e(al_ccabc055[8]),
    .f(al_7b4ebd2a),
    .o(al_2418b5af));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_7f0b20e (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_2418b5af),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[8]),
    .f(al_b24d99c7[7]),
    .o(al_bde0dc95[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h084c2a6e195d3b7f))
    al_265c026d (
    .a(al_8db3355a),
    .b(al_dd37dc5d),
    .c(al_35d85285[7]),
    .d(al_46ea2d9f[9]),
    .e(al_ccabc055[9]),
    .f(al_e3fa27d),
    .o(al_4a696460));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*~(C)*~(A)+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*~(A)+~(~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B)))*C*A+~(E*~(F)*~((D*B))+E*F*~((D*B))+~(E)*F*(D*B)+E*F*(D*B))*C*A)"),
    .INIT(64'h5f5f4e0a1b5f0a0a))
    al_fb9cd108 (
    .a(al_6f809586),
    .b(al_e87ca79),
    .c(al_4a696460),
    .d(al_3f1d46e5),
    .e(al_a16ef20a[9]),
    .f(al_b24d99c7[8]),
    .o(al_bde0dc95[9]));
  AL_DFF_X al_8034d3e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e2d7fc47),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f56de171));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_c260bdd2 (
    .a(al_fccc3291),
    .b(al_9c16c2f5),
    .c(al_126b3afd[1]),
    .o(al_d485b6de));
  AL_MAP_LUT5 #(
    .EQN("(A*(B*~(C)*D*~(E)+~(B)*~(C)*~(D)*E+~(B)*C*~(D)*E+~(B)*~(C)*D*E+B*~(C)*D*E+~(B)*C*D*E+B*C*D*E))"),
    .INIT(32'haa220800))
    al_d5dba9b8 (
    .a(al_b8437eb4),
    .b(al_1d3bfd2e),
    .c(al_d485b6de),
    .d(al_d72f4570),
    .e(al_bccf82af),
    .o(al_e72a5b80));
  AL_DFF_X al_1f9b0784 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e72a5b80),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bccf82af));
  AL_DFF_X al_ac11802 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0b8db17),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a2250ee));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~C*B*~(~E*~D)))"),
    .INIT(32'ha2a2a2aa))
    al_d892d215 (
    .a(al_1d3bfd2e),
    .b(al_d72f4570),
    .c(al_bccf82af),
    .d(al_9c16c2f5),
    .e(al_126b3afd[1]),
    .o(al_2d6e7982));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    al_38f5f0ba (
    .a(al_2d6e7982),
    .b(al_b8437eb4),
    .c(al_37a2cec8),
    .d(al_9c16c2f5),
    .o(al_61085a1a));
  AL_DFF_X al_ca77ef82 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_61085a1a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c16c2f5));
  AL_DFF_X al_c4ccf2a1 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(1'b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0ecd262));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_b4dd8101 (
    .a(al_6a0e908c),
    .b(al_2c3e73df),
    .o(al_fa66b6a3));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*C*~A))"),
    .INIT(16'hdccc))
    al_c3dcbe9b (
    .a(al_a25a6119),
    .b(al_cc4ef047),
    .c(al_fa66b6a3),
    .d(al_519869c),
    .o(al_536fd7fd));
  AL_DFF_X al_3549c766 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_536fd7fd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_519869c));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_8f08b457 (
    .a(1'b0),
    .o({al_24cba21e,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_495af386 (
    .a(al_126b3afd[2]),
    .b(al_519869c),
    .c(al_24cba21e),
    .o({al_6cfd8dcf,al_683f5875[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2d64e6b8 (
    .a(al_126b3afd[3]),
    .b(1'b0),
    .c(al_6cfd8dcf),
    .o({al_a2aa312d,al_683f5875[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_82d0e41c (
    .a(al_126b3afd[4]),
    .b(1'b0),
    .c(al_a2aa312d),
    .o({al_5beecaa3,al_683f5875[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d373e6a4 (
    .a(al_126b3afd[5]),
    .b(1'b0),
    .c(al_5beecaa3),
    .o({al_3b6c54b6,al_683f5875[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f3e4fc09 (
    .a(al_126b3afd[6]),
    .b(1'b0),
    .c(al_3b6c54b6),
    .o({al_50439dee,al_683f5875[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d3598443 (
    .a(al_126b3afd[7]),
    .b(1'b0),
    .c(al_50439dee),
    .o({al_72de3c0a,al_683f5875[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_db91bc2b (
    .a(al_126b3afd[8]),
    .b(1'b0),
    .c(al_72de3c0a),
    .o({al_b0555243,al_683f5875[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5416914a (
    .a(al_126b3afd[9]),
    .b(1'b0),
    .c(al_b0555243),
    .o({al_210b38e6,al_683f5875[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a98e6772 (
    .a(al_126b3afd[10]),
    .b(1'b0),
    .c(al_210b38e6),
    .o({al_bbee20b8,al_683f5875[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_59dc3e92 (
    .a(al_126b3afd[11]),
    .b(1'b0),
    .c(al_bbee20b8),
    .o({al_c1d3ffb3,al_683f5875[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5690057a (
    .a(al_126b3afd[12]),
    .b(1'b0),
    .c(al_c1d3ffb3),
    .o({al_3e1875be,al_683f5875[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f9041b78 (
    .a(al_126b3afd[13]),
    .b(1'b0),
    .c(al_3e1875be),
    .o({al_27878642,al_683f5875[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_52a8cbfe (
    .a(al_126b3afd[14]),
    .b(1'b0),
    .c(al_27878642),
    .o({al_ac867fa2,al_683f5875[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3874dbfd (
    .a(al_126b3afd[15]),
    .b(1'b0),
    .c(al_ac867fa2),
    .o({al_8b9b5b1d,al_683f5875[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_64fd65d (
    .a(al_126b3afd[16]),
    .b(1'b0),
    .c(al_8b9b5b1d),
    .o({al_80a6299b,al_683f5875[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a420e51e (
    .a(al_126b3afd[17]),
    .b(1'b0),
    .c(al_80a6299b),
    .o({al_6305766,al_683f5875[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_926c3cd0 (
    .a(al_126b3afd[18]),
    .b(1'b0),
    .c(al_6305766),
    .o({al_e51dc3c,al_683f5875[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9d2987c (
    .a(al_126b3afd[19]),
    .b(1'b0),
    .c(al_e51dc3c),
    .o({al_5fe5e97d,al_683f5875[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a5288bde (
    .a(al_126b3afd[20]),
    .b(1'b0),
    .c(al_5fe5e97d),
    .o({al_35379d79,al_683f5875[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_479aaabb (
    .a(al_126b3afd[21]),
    .b(1'b0),
    .c(al_35379d79),
    .o({al_5a3ca2c7,al_683f5875[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_755fe1ba (
    .a(al_126b3afd[22]),
    .b(1'b0),
    .c(al_5a3ca2c7),
    .o({al_e791df33,al_683f5875[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c6e4649c (
    .a(al_126b3afd[23]),
    .b(1'b0),
    .c(al_e791df33),
    .o({al_168ce6c3,al_683f5875[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9f62d15c (
    .a(al_126b3afd[24]),
    .b(1'b0),
    .c(al_168ce6c3),
    .o({al_1e8c20b0,al_683f5875[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d1d31b29 (
    .a(al_126b3afd[25]),
    .b(1'b0),
    .c(al_1e8c20b0),
    .o({al_5a6794e3,al_683f5875[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_22ccd57 (
    .a(al_126b3afd[26]),
    .b(1'b0),
    .c(al_5a6794e3),
    .o({al_d3114685,al_683f5875[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a276e1ab (
    .a(al_126b3afd[27]),
    .b(1'b0),
    .c(al_d3114685),
    .o({al_4ea1bb54,al_683f5875[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3e377cf0 (
    .a(al_126b3afd[28]),
    .b(1'b0),
    .c(al_4ea1bb54),
    .o({al_d5e048cf,al_683f5875[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_58385790 (
    .a(al_126b3afd[29]),
    .b(1'b0),
    .c(al_d5e048cf),
    .o({al_1eaad5d4,al_683f5875[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4731f73 (
    .a(al_126b3afd[30]),
    .b(1'b0),
    .c(al_1eaad5d4),
    .o({al_c63ed4c6,al_683f5875[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f7b4626d (
    .a(al_126b3afd[31]),
    .b(1'b0),
    .c(al_c63ed4c6),
    .o({open_n11,al_683f5875[29]}));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_9444382f (
    .a(al_4ed450cb),
    .b(al_fa66b6a3),
    .c(al_683f5875[8]),
    .o(al_c1211126[10]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_35dc14be (
    .a(al_667db93d),
    .b(al_fa66b6a3),
    .c(al_683f5875[9]),
    .o(al_c1211126[11]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_e986bf6e (
    .a(al_fb26226a),
    .b(al_fa66b6a3),
    .c(al_683f5875[10]),
    .o(al_c1211126[12]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_9219de58 (
    .a(al_c4d4b7f5),
    .b(al_fa66b6a3),
    .c(al_683f5875[11]),
    .o(al_c1211126[13]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_a20eac6a (
    .a(al_13708b94),
    .b(al_fa66b6a3),
    .c(al_683f5875[12]),
    .o(al_c1211126[14]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_4678a7b6 (
    .a(al_8cb8f5f5),
    .b(al_fa66b6a3),
    .c(al_683f5875[13]),
    .o(al_c1211126[15]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_7dfa4907 (
    .a(al_c5cc2f9b),
    .b(al_fa66b6a3),
    .c(al_683f5875[14]),
    .o(al_c1211126[16]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_8a7d5392 (
    .a(al_c048f5a0),
    .b(al_fa66b6a3),
    .c(al_683f5875[15]),
    .o(al_c1211126[17]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_9ae2cd2d (
    .a(al_c6cd8be8),
    .b(al_fa66b6a3),
    .c(al_683f5875[16]),
    .o(al_c1211126[18]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_2184de51 (
    .a(al_31822056),
    .b(al_fa66b6a3),
    .c(al_683f5875[17]),
    .o(al_c1211126[19]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D*~C*B))"),
    .INIT(16'h5d55))
    al_cde62e11 (
    .a(al_81e43d4),
    .b(al_fa66b6a3),
    .c(al_519869c),
    .d(al_126b3afd[1]),
    .o(al_c1211126[1]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_383623e2 (
    .a(al_6e8dae0d),
    .b(al_fa66b6a3),
    .c(al_683f5875[18]),
    .o(al_c1211126[20]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_3c6a6302 (
    .a(al_f76f8d54),
    .b(al_fa66b6a3),
    .c(al_683f5875[19]),
    .o(al_c1211126[21]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_730b74d2 (
    .a(al_825438f5),
    .b(al_fa66b6a3),
    .c(al_683f5875[20]),
    .o(al_c1211126[22]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_ca2df481 (
    .a(al_ab46d2b9),
    .b(al_fa66b6a3),
    .c(al_683f5875[21]),
    .o(al_c1211126[23]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_f9b2cd6e (
    .a(al_d33dd538),
    .b(al_fa66b6a3),
    .c(al_683f5875[22]),
    .o(al_c1211126[24]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_d4ef67f7 (
    .a(al_b62de081),
    .b(al_fa66b6a3),
    .c(al_683f5875[23]),
    .o(al_c1211126[25]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_28186e6f (
    .a(al_447f0158),
    .b(al_fa66b6a3),
    .c(al_683f5875[24]),
    .o(al_c1211126[26]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_f3208bed (
    .a(al_a0670bff),
    .b(al_fa66b6a3),
    .c(al_683f5875[25]),
    .o(al_c1211126[27]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_3a515181 (
    .a(al_74973e72),
    .b(al_fa66b6a3),
    .c(al_683f5875[26]),
    .o(al_c1211126[28]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_d0f7155b (
    .a(al_cae3c642),
    .b(al_fa66b6a3),
    .c(al_683f5875[27]),
    .o(al_c1211126[29]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_5764139f (
    .a(al_3db1ed2d),
    .b(al_fa66b6a3),
    .c(al_683f5875[0]),
    .o(al_c1211126[2]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_f6a827b0 (
    .a(al_ac5b8836),
    .b(al_fa66b6a3),
    .c(al_683f5875[28]),
    .o(al_c1211126[30]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_554ebdec (
    .a(al_9bb19ed8),
    .b(al_fa66b6a3),
    .c(al_683f5875[29]),
    .o(al_c1211126[31]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_818428c4 (
    .a(al_e9dadc09),
    .b(al_fa66b6a3),
    .c(al_683f5875[1]),
    .o(al_c1211126[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_86e1af1b (
    .a(al_3be09bce),
    .b(al_fa66b6a3),
    .c(al_683f5875[2]),
    .o(al_c1211126[4]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_704eb298 (
    .a(al_8773b31),
    .b(al_fa66b6a3),
    .c(al_683f5875[3]),
    .o(al_c1211126[5]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_ceeee03f (
    .a(al_640ea1c6),
    .b(al_fa66b6a3),
    .c(al_683f5875[4]),
    .o(al_c1211126[6]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_7dcc3625 (
    .a(al_4e819ed5),
    .b(al_fa66b6a3),
    .c(al_683f5875[5]),
    .o(al_c1211126[7]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_4d523a44 (
    .a(al_2418b5af),
    .b(al_fa66b6a3),
    .c(al_683f5875[6]),
    .o(al_c1211126[8]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_ce910ace (
    .a(al_4a696460),
    .b(al_fa66b6a3),
    .c(al_683f5875[7]),
    .o(al_c1211126[9]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_2fb5e708 (
    .i(al_a16ef20a[0]),
    .o(al_adeed2de[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_97cdc33 (
    .i(al_adeed2de[0]),
    .o(al_4d016a39));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f455a80f (
    .i(al_8d9bdfff),
    .o(al_adeed2de[10]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_ecaa2272 (
    .i(al_adeed2de[10]),
    .o(al_2cd19c12));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_cd53b264 (
    .i(al_70f172be),
    .o(al_adeed2de[11]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_21819ee (
    .i(al_adeed2de[11]),
    .o(al_cc989ac9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_51ac9685 (
    .i(al_c89d1229),
    .o(al_adeed2de[12]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9955da60 (
    .i(al_adeed2de[12]),
    .o(al_1953385a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4c815fc4 (
    .i(al_2d354b),
    .o(al_adeed2de[13]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6fb741ca (
    .i(al_adeed2de[13]),
    .o(al_be6e0599));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c1b50741 (
    .i(al_2fb7633),
    .o(al_adeed2de[14]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1fc80884 (
    .i(al_adeed2de[14]),
    .o(al_afe5948f));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8f35a715 (
    .i(al_5b3ba944),
    .o(al_adeed2de[15]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3dab82b (
    .i(al_adeed2de[15]),
    .o(al_d1fc8906));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_24393d1d (
    .i(al_f5f3edb6),
    .o(al_adeed2de[16]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d3c5c9db (
    .i(al_adeed2de[16]),
    .o(al_9df5b848));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_894a1aea (
    .i(al_d0702be9),
    .o(al_adeed2de[17]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d8b706e8 (
    .i(al_adeed2de[17]),
    .o(al_afd990ff));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f0b7d598 (
    .i(al_2eb5050b),
    .o(al_adeed2de[18]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_492ce43e (
    .i(al_adeed2de[18]),
    .o(al_7bf844c2));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_84896047 (
    .i(al_89a93b84),
    .o(al_adeed2de[19]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_5fa37784 (
    .i(al_adeed2de[19]),
    .o(al_b6803a27));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3b263fc4 (
    .i(al_e79b3dfa),
    .o(al_adeed2de[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b53fdfa6 (
    .i(al_adeed2de[1]),
    .o(al_6ae2a07d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_471e3543 (
    .i(al_82b168eb),
    .o(al_adeed2de[20]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_aa515187 (
    .i(al_adeed2de[20]),
    .o(al_20b06ef3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3d6b3e4d (
    .i(al_e2259475),
    .o(al_adeed2de[21]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e46b0eac (
    .i(al_adeed2de[21]),
    .o(al_b40171bd));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_16ef8343 (
    .i(al_6758eae2),
    .o(al_adeed2de[22]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_758c26f2 (
    .i(al_adeed2de[22]),
    .o(al_42b103ed));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_34a3f8e4 (
    .i(al_f814979a),
    .o(al_adeed2de[23]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4bd1f87d (
    .i(al_adeed2de[23]),
    .o(al_5a93aea7));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4c1dc222 (
    .i(al_5ca98598),
    .o(al_adeed2de[24]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_bca3445f (
    .i(al_adeed2de[24]),
    .o(al_40d63aa3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7a4fc84c (
    .i(al_267d2aa),
    .o(al_adeed2de[25]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_f281ff3e (
    .i(al_adeed2de[25]),
    .o(al_89782fa0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_9aaaea3f (
    .i(al_debfa536),
    .o(al_adeed2de[26]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_df998b0 (
    .i(al_adeed2de[26]),
    .o(al_faaecf2));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8b64186b (
    .i(al_f19f190e),
    .o(al_adeed2de[27]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_51ee8acb (
    .i(al_adeed2de[27]),
    .o(al_ad2a00e5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_43e09905 (
    .i(al_9852e0df),
    .o(al_adeed2de[28]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_f7f38e4d (
    .i(al_adeed2de[28]),
    .o(al_193c583f));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_9909def5 (
    .i(al_ecd761fc),
    .o(al_adeed2de[29]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_bbf5f3bf (
    .i(al_adeed2de[29]),
    .o(al_a155e0b3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a79347a6 (
    .i(al_ca581e6c),
    .o(al_adeed2de[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_459e4cce (
    .i(al_adeed2de[2]),
    .o(al_cc5bfca5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_920f922 (
    .i(al_c64cf9f6),
    .o(al_adeed2de[30]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_840a98d2 (
    .i(al_adeed2de[30]),
    .o(al_89bb053a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_413e5d96 (
    .i(al_5e07bd5e),
    .o(al_adeed2de[31]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_5199781a (
    .i(al_adeed2de[31]),
    .o(al_4efe0c98));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c4afae62 (
    .i(al_428b50b6),
    .o(al_adeed2de[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1bf673b4 (
    .i(al_adeed2de[3]),
    .o(al_5bcd7a0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_6fab13a1 (
    .i(al_a3f3ee06),
    .o(al_adeed2de[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e58c6ddc (
    .i(al_adeed2de[4]),
    .o(al_3ab03292));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5f41dc7 (
    .i(al_263322e4),
    .o(al_adeed2de[5]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_5459ff91 (
    .i(al_adeed2de[5]),
    .o(al_22da7862));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_6f45535b (
    .i(al_63bbd3a2),
    .o(al_adeed2de[6]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_421f3a2a (
    .i(al_adeed2de[6]),
    .o(al_45322fba));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5a639723 (
    .i(al_6ab73d4d),
    .o(al_adeed2de[7]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c63b8674 (
    .i(al_adeed2de[7]),
    .o(al_c585508d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7727b20b (
    .i(al_fd8d8e0c),
    .o(al_adeed2de[8]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3caa25a9 (
    .i(al_adeed2de[8]),
    .o(al_7b4ebd2a));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_51f84a2 (
    .i(al_a89113a9),
    .o(al_adeed2de[9]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_895edc87 (
    .i(al_adeed2de[9]),
    .o(al_e3fa27d));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*A))+D*C*~((~B*A))+~(D)*C*(~B*A)+D*C*(~B*A))"),
    .INIT(16'hfd20))
    al_2366ba43 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[19]),
    .d(al_85a2bdb0[31]),
    .o(al_8c22c3eb));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*A))+D*C*~((~B*A))+~(D)*C*(~B*A)+D*C*(~B*A))"),
    .INIT(16'hfd20))
    al_4dfb8835 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[18]),
    .d(al_85a2bdb0[31]),
    .o(al_cc14dad7));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*A))+D*C*~((~B*A))+~(D)*C*(~B*A)+D*C*(~B*A))"),
    .INIT(16'hfd20))
    al_c673e072 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[17]),
    .d(al_85a2bdb0[31]),
    .o(al_4bfb7d3a));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*A))+D*C*~((~B*A))+~(D)*C*(~B*A)+D*C*(~B*A))"),
    .INIT(16'hfd20))
    al_f3626ae1 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[16]),
    .d(al_85a2bdb0[31]),
    .o(al_bcf22cd5));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*A))+D*C*~((~B*A))+~(D)*C*(~B*A)+D*C*(~B*A))"),
    .INIT(16'hfd20))
    al_225fb924 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[15]),
    .d(al_85a2bdb0[31]),
    .o(al_96c3cafb));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*A))+D*C*~((~B*A))+~(D)*C*(~B*A)+D*C*(~B*A))"),
    .INIT(16'hfd20))
    al_93aa55fb (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[14]),
    .d(al_85a2bdb0[31]),
    .o(al_2cce4860));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*A))+D*C*~((~B*A))+~(D)*C*(~B*A)+D*C*(~B*A))"),
    .INIT(16'hfd20))
    al_bb0a73d3 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[13]),
    .d(al_85a2bdb0[31]),
    .o(al_420d5318));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*A))+D*C*~((~B*A))+~(D)*C*(~B*A)+D*C*(~B*A))"),
    .INIT(16'hfd20))
    al_b7beba87 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[12]),
    .d(al_85a2bdb0[31]),
    .o(al_383f9835));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*A))+C*D*~((~B*A))+~(C)*D*(~B*A)+C*D*(~B*A))"),
    .INIT(16'hf2d0))
    al_27ce8e4f (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[7]),
    .d(al_85a2bdb0[20]),
    .o(al_1405651f));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*A))+C*D*~((~B*A))+~(C)*D*(~B*A)+C*D*(~B*A))"),
    .INIT(16'hf2d0))
    al_91d7928b (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[11]),
    .d(al_85a2bdb0[24]),
    .o(al_a40c439));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*A))+C*D*~((~B*A))+~(C)*D*(~B*A)+C*D*(~B*A))"),
    .INIT(16'hf2d0))
    al_f32a8f9 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[10]),
    .d(al_85a2bdb0[23]),
    .o(al_de666865));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*A))+C*D*~((~B*A))+~(C)*D*(~B*A)+C*D*(~B*A))"),
    .INIT(16'hf2d0))
    al_e32c3195 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[9]),
    .d(al_85a2bdb0[22]),
    .o(al_4cc97ac1));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*A))+C*D*~((~B*A))+~(C)*D*(~B*A)+C*D*(~B*A))"),
    .INIT(16'hf2d0))
    al_4465bad0 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[8]),
    .d(al_85a2bdb0[21]),
    .o(al_1d7074bf));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_de7c8918 (
    .a(al_acd38e8e),
    .b(al_d518b626),
    .o(al_4736f54a));
  AL_DFF_X al_bffe421c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[7]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[8]));
  AL_DFF_X al_2b03af3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[8]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[9]));
  AL_DFF_X al_1edfc532 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[9]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[10]));
  AL_DFF_X al_67df7702 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[10]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[11]));
  AL_DFF_X al_8aa6b08e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[11]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[12]));
  AL_DFF_X al_efb17dfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[12]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[13]));
  AL_DFF_X al_aaca23ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[13]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[14]));
  AL_DFF_X al_9db78a12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[14]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[15]));
  AL_DFF_X al_93af0048 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[15]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[16]));
  AL_DFF_X al_46abb091 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[16]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[17]));
  AL_DFF_X al_f458b215 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRESP),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[0]));
  AL_DFF_X al_4b665528 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[17]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[18]));
  AL_DFF_X al_4cb3e186 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[18]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[19]));
  AL_DFF_X al_7e40bfe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[19]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[20]));
  AL_DFF_X al_6012d2d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[20]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[21]));
  AL_DFF_X al_345f1431 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[21]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[22]));
  AL_DFF_X al_4131fc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[22]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[23]));
  AL_DFF_X al_bdb0e467 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[23]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[24]));
  AL_DFF_X al_194d260d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[24]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[25]));
  AL_DFF_X al_d5a7178 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[25]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[26]));
  AL_DFF_X al_508ad212 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[26]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[27]));
  AL_DFF_X al_1439a22c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[0]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[1]));
  AL_DFF_X al_f3b4b157 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[27]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[28]));
  AL_DFF_X al_1c0e4604 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[28]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[29]));
  AL_DFF_X al_cb62a13c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[29]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[30]));
  AL_DFF_X al_d7a00e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[30]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[31]));
  AL_DFF_X al_71b1ed59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[31]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[32]));
  AL_DFF_X al_544d4cac (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[1]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[2]));
  AL_DFF_X al_11b74881 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[2]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[3]));
  AL_DFF_X al_759dea3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[3]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[4]));
  AL_DFF_X al_2b17de10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[4]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[5]));
  AL_DFF_X al_af671c5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[5]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[6]));
  AL_DFF_X al_289538e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(iBusAhb_HRDATA[6]),
    .en(al_4736f54a),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b86dd14b[7]));
  AL_DFF_X al_6604197 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2b6037c7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d518b626));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9375b36e (
    .a(al_523a156f),
    .b(al_e0005a94),
    .o(al_2b6037c7));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h4c194613))
    al_6afb6d98 (
    .a(al_b8437eb4),
    .b(al_e0005a94),
    .c(al_7a486383),
    .d(al_9b5530fd[0]),
    .e(al_202f2c67[0]),
    .o(al_b537d840[0]));
  AL_MAP_LUT4 #(
    .EQN("(~((~B*~A))*~(C)*~(D)+(~B*~A)*~(C)*~(D)+(~B*~A)*C*~(D)+~((~B*~A))*~(C)*D+(~B*~A)*C*D)"),
    .INIT(16'h1e1f))
    al_d52f8373 (
    .a(al_e0005a94),
    .b(al_202f2c67[0]),
    .c(al_202f2c67[1]),
    .d(al_202f2c67[2]),
    .o(al_b2f6a2a2));
  AL_MAP_LUT4 #(
    .EQN("~(~(D@A)*~(C)*~(B)+~(D@A)*C*~(B)+~(~(D@A))*C*B+~(D@A)*C*B)"),
    .INIT(16'h1d2e))
    al_2acc9d06 (
    .a(al_cd3394ba),
    .b(al_b8437eb4),
    .c(al_b2f6a2a2),
    .d(al_9b5530fd[1]),
    .o(al_b537d840[1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_4af8f31 (
    .a(al_c795a432),
    .b(al_a8151162),
    .c(al_2c3e73df),
    .o(al_b8437eb4));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_d316dea2 (
    .a(al_e0005a94),
    .b(al_9b5530fd[0]),
    .o(al_cd3394ba));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    al_95d334ad (
    .a(al_e0005a94),
    .b(al_202f2c67[0]),
    .c(al_202f2c67[1]),
    .d(al_202f2c67[2]),
    .o(al_2978b178[2]));
  AL_MAP_LUT5 #(
    .EQN("((E@(~D*A))*~(C)*~(B)+(E@(~D*A))*C*~(B)+~((E@(~D*A)))*C*B+(E@(~D*A))*C*B)"),
    .INIT(32'hf3d1c0e2))
    al_456842f7 (
    .a(al_cd3394ba),
    .b(al_b8437eb4),
    .c(al_2978b178[2]),
    .d(al_9b5530fd[1]),
    .e(al_9b5530fd[2]),
    .o(al_b537d840[2]));
  AL_DFF_X al_515ac502 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(1'b0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d334d88));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    al_e1538c93 (
    .a(al_3f1d46e5),
    .b(al_a7b01c14[2]),
    .c(al_f6cd735f),
    .d(al_69807e37),
    .o(al_fa0903ac));
  AL_DFF_X al_1ec5f5fc (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_fa0903ac),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a2deaa78));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_c06487d (
    .a(al_24a3e858),
    .o(al_6515336d[2]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*B*~(~D*C)))"),
    .INIT(32'heeaeaaaa))
    al_2e810bc8 (
    .a(al_cc4ef047),
    .b(al_b8437eb4),
    .c(al_1d3bfd2e),
    .d(al_37a2cec8),
    .e(al_f49992c3),
    .o(al_94c23c7d));
  AL_DFF_X al_c9e4eb95 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_94c23c7d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f49992c3));
  AL_DFF_X al_fd27a9d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f14f6e5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24a3e858));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_498a805f (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_24a3e858),
    .o(al_6f14f6e5));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_f3bc540d (
    .a(al_85a2bdb0[12]),
    .o(al_b63bb946));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~A*~(D*~B)))*~(C)+~E*(~A*~(D*~B))*~(C)+~(~E)*(~A*~(D*~B))*C+~E*(~A*~(D*~B))*C)"),
    .INIT(32'hbfafb0a0))
    al_d5bb3554 (
    .a(al_2a0680fd),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[0]),
    .e(al_25fbce42[32]),
    .o(al_1f3eaa15[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6ffd740a (
    .a(iBusAhb_HRDATA[26]),
    .b(al_b86dd14b[27]),
    .c(al_d518b626),
    .o(al_cf18c1c6[26]));
  AL_MAP_LUT6 #(
    .EQN("(F*~((E*~((~C*~A))*~(B)+E*(~C*~A)*~(B)+~(E)*(~C*~A)*B+E*(~C*~A)*B))*~(D)+F*(E*~((~C*~A))*~(B)+E*(~C*~A)*~(B)+~(E)*(~C*~A)*B+E*(~C*~A)*B)*~(D)+~(F)*(E*~((~C*~A))*~(B)+E*(~C*~A)*~(B)+~(E)*(~C*~A)*B+E*(~C*~A)*B)*D+F*(E*~((~C*~A))*~(B)+E*(~C*~A)*~(B)+~(E)*(~C*~A)*B+E*(~C*~A)*B)*D)"),
    .INIT(64'h37ff04ff37000400))
    al_c3759ac7 (
    .a(al_6e7063d6),
    .b(al_a7b01c14[2]),
    .c(al_8647937a),
    .d(al_8905c135),
    .e(al_85a2bdb0[10]),
    .f(al_25fbce42[42]),
    .o(al_1f3eaa15[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2441cdfb (
    .a(iBusAhb_HRDATA[10]),
    .b(al_b86dd14b[11]),
    .c(al_d518b626),
    .o(al_cf18c1c6[10]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_b115f71 (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[26]),
    .c(al_cf18c1c6[10]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_d344e0e5));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_fb56fa38 (
    .a(al_d344e0e5),
    .b(al_e2d7fc47),
    .c(al_5fd02584[10]),
    .o(al_2d35601b));
  AL_MAP_LUT6 #(
    .EQN("(~B*(~(A)*C*~(D)*~(E)*~(F)+A*C*~(D)*~(E)*~(F)+~(A)*C*D*~(E)*~(F)+A*C*D*~(E)*~(F)+~(A)*~(C)*~(D)*E*~(F)+A*~(C)*~(D)*E*~(F)+~(A)*C*~(D)*E*~(F)+A*C*~(D)*E*~(F)+~(A)*~(C)*D*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*D*E*~(F)+~(A)*~(C)*~(D)*E*F+A*~(C)*~(D)*E*F+A*C*~(D)*E*F))"),
    .INIT(64'h0023000033333030))
    al_2ae43e45 (
    .a(al_955e8db5),
    .b(al_4002af45),
    .c(al_843f038d),
    .d(al_ba3f2ea7),
    .e(al_7a7cc81),
    .f(al_2d35601b),
    .o(al_6e7063d6));
  AL_MAP_LUT6 #(
    .EQN("(A*~(C)*~((~D*~B))*~(E)*~(F)+~(A)*C*~((~D*~B))*~(E)*~(F)+A*C*~((~D*~B))*~(E)*~(F)+A*~(C)*(~D*~B)*~(E)*~(F)+~(A)*C*(~D*~B)*~(E)*~(F)+A*C*(~D*~B)*~(E)*~(F)+A*~(C)*~((~D*~B))*E*~(F)+~(A)*C*~((~D*~B))*E*~(F)+A*C*~((~D*~B))*E*~(F)+~(A)*C*(~D*~B)*E*~(F)+A*C*(~D*~B)*E*~(F)+~(A)*C*~((~D*~B))*~(E)*F+~(A)*C*(~D*~B)*~(E)*F+A*C*(~D*~B)*~(E)*F+~(A)*C*~((~D*~B))*E*F+~(A)*C*(~D*~B)*E*F+A*C*(~D*~B)*E*F)"),
    .INIT(64'h50705070faf8fafa))
    al_fdadf9e6 (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_1f0371f8),
    .d(al_ba3f2ea7),
    .e(al_7a7cc81),
    .f(al_2d35601b),
    .o(al_8647937a));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_64bd98e6 (
    .a(iBusAhb_HRDATA[27]),
    .b(al_b86dd14b[28]),
    .c(al_d518b626),
    .o(al_cf18c1c6[27]));
  AL_MAP_LUT5 #(
    .EQN("(E*~((D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))*~(C)+E*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*~(C)+~(E)*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C+E*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C)"),
    .INIT(32'hbf8fb080))
    al_eedad5ce (
    .a(al_8778492e[11]),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[11]),
    .e(al_25fbce42[43]),
    .o(al_1f3eaa15[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_af948b45 (
    .a(iBusAhb_HRDATA[11]),
    .b(al_b86dd14b[12]),
    .c(al_d518b626),
    .o(al_cf18c1c6[11]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_b97d1edf (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[27]),
    .c(al_cf18c1c6[11]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_87b30ed5));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_2839ec06 (
    .a(al_87b30ed5),
    .b(al_e2d7fc47),
    .c(al_5fd02584[11]),
    .o(al_e22f5efa));
  AL_MAP_LUT6 #(
    .EQN("(F*(~(A)*~(C)*~((~D*~B))*~(E)+A*~(C)*~((~D*~B))*~(E)+A*C*~((~D*~B))*~(E)+~(A)*~(C)*(~D*~B)*~(E)+A*~(C)*(~D*~B)*~(E)+~(A)*~(C)*~((~D*~B))*E+A*~(C)*~((~D*~B))*E+A*C*~((~D*~B))*E))"),
    .INIT(64'haf8caf8f00000000))
    al_b9b49093 (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_1f0371f8),
    .d(al_ba3f2ea7),
    .e(al_7a7cc81),
    .f(al_e22f5efa),
    .o(al_286b6a5c));
  AL_MAP_LUT6 #(
    .EQN("(A*~(~C*(~D*~((~E*B))*~(F)+~D*(~E*B)*~(F)+~(~D)*(~E*B)*F+~D*(~E*B)*F)))"),
    .INIT(64'haaaaa2a2aaa0aaa0))
    al_ba3a72f5 (
    .a(al_286b6a5c),
    .b(al_955e8db5),
    .c(al_4002af45),
    .d(al_843f038d),
    .e(al_ba3f2ea7),
    .f(al_7a7cc81),
    .o(al_8778492e[11]));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(F*E*~(D*C)))"),
    .INIT(64'h8000888888888888))
    al_aab087ff (
    .a(al_c7467d2d),
    .b(al_7a7cc81),
    .c(al_55bbd6fb),
    .d(al_8f175a04),
    .e(al_2d35601b),
    .f(al_e22f5efa),
    .o(al_74e1f810));
  AL_MAP_LUT6 #(
    .EQN("(B*~(~E*~((~D*~(F*~A)))*~(C)+~E*(~D*~(F*~A))*~(C)+~(~E)*(~D*~(F*~A))*C+~E*(~D*~(F*~A))*C))"),
    .INIT(64'hcc4cc040cc0cc000))
    al_c62ce9f9 (
    .a(al_90d6c009),
    .b(al_1f0371f8),
    .c(al_ba3f2ea7),
    .d(al_7a7cc81),
    .e(al_3f6865d3),
    .f(al_78e2749c),
    .o(al_5c743358));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_738706d9 (
    .a(al_e1adfd34),
    .b(al_ba3f2ea7),
    .c(al_7a7cc81),
    .o(al_f4b0c1c2[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(C)*~((~D*~B))*~(E)*~(F)+~(A)*~(C)*~((~D*~B))*E*~(F)+A*~(C)*~((~D*~B))*E*~(F)+A*~(C)*(~D*~B)*E*~(F)+~(A)*~(C)*~((~D*~B))*~(E)*F+~(A)*~(C)*~((~D*~B))*E*F+A*~(C)*~((~D*~B))*E*F+~(A)*C*~((~D*~B))*E*F+A*C*~((~D*~B))*E*F+A*~(C)*(~D*~B)*E*F+~(A)*C*(~D*~B)*E*F+A*C*(~D*~B)*E*F)"),
    .INIT(64'hfffe05040f0e0504))
    al_56983355 (
    .a(al_74e1f810),
    .b(al_5c743358),
    .c(al_bdf9a7dd),
    .d(al_f4b0c1c2[12]),
    .e(al_4002af45),
    .f(al_3f6865d3),
    .o(al_8778492e[12]));
  AL_MAP_LUT5 #(
    .EQN("(E*~((D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))*~(C)+E*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*~(C)+~(E)*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C+E*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C)"),
    .INIT(32'hbf8fb080))
    al_3ac24f64 (
    .a(al_8778492e[12]),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[12]),
    .e(al_25fbce42[44]),
    .o(al_1f3eaa15[12]));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(F*~((~E*C*~A))*~(D)+F*(~E*C*~A)*~(D)+~(F)*(~E*C*~A)*D+F*(~E*C*~A)*D))"),
    .INIT(64'h3300230033332333))
    al_880fb104 (
    .a(al_90d6c009),
    .b(al_843f038d),
    .c(al_f65e6902[3]),
    .d(al_ba3f2ea7),
    .e(al_7a7cc81),
    .f(al_3f6865d3),
    .o(al_6df79c7b));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*~B))"),
    .INIT(16'h4500))
    al_fa71d206 (
    .a(al_843f038d),
    .b(al_55bbd6fb),
    .c(al_2d35601b),
    .d(al_e22f5efa),
    .o(al_7c75aadd));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(C)*~(D)*~(E)*~((F*B))+A*~(C)*~(D)*~(E)*~((F*B))+~(A)*C*~(D)*~(E)*~((F*B))+A*C*~(D)*~(E)*~((F*B))+~(A)*~(C)*D*~(E)*~((F*B))+A*~(C)*D*~(E)*~((F*B))+A*C*D*~(E)*~((F*B))+~(A)*C*~(D)*E*~((F*B))+A*C*~(D)*E*~((F*B))+~(A)*~(C)*D*E*~((F*B))+A*~(C)*D*E*~((F*B))+A*C*D*E*~((F*B))+~(A)*~(C)*~(D)*~(E)*(F*B)+A*~(C)*~(D)*~(E)*(F*B)+~(A)*~(C)*D*~(E)*(F*B)+A*~(C)*D*~(E)*(F*B)+A*C*D*~(E)*(F*B)+~(A)*C*~(D)*E*(F*B)+A*C*~(D)*E*(F*B)+~(A)*~(C)*D*E*(F*B)+A*~(C)*D*E*(F*B)+A*C*D*E*(F*B))"),
    .INIT(64'haff0af3faff0afff))
    al_9aeee76c (
    .a(al_6df79c7b),
    .b(al_7c75aadd),
    .c(al_4002af45),
    .d(al_1f0371f8),
    .e(al_ba3f2ea7),
    .f(al_7a7cc81),
    .o(al_f7b11965));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B))*~(C)+~E*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*~(C)+~(~E)*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*C+~E*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*C)"),
    .INIT(32'h7f4f7040))
    al_8330cc76 (
    .a(al_f7b11965),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[13]),
    .e(al_25fbce42[45]),
    .o(al_1f3eaa15[13]));
  AL_MAP_LUT5 #(
    .EQN("(~C*~A*~(E*D*~B))"),
    .INIT(32'h04050505))
    al_849b8b81 (
    .a(al_7c8ae043),
    .b(al_bd10bda8),
    .c(al_1f0371f8),
    .d(al_2d35601b),
    .e(al_e22f5efa),
    .o(al_83a071a4));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(C*~(~(E*~D)*~(F*A))))"),
    .INIT(64'h1303131333033333))
    al_9d8d5327 (
    .a(al_73767b69),
    .b(al_83a071a4),
    .c(al_1f0371f8),
    .d(al_ba3f2ea7),
    .e(al_3f6865d3),
    .f(al_f65e6902[4]),
    .o(al_55ed4df1));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_9be46749 (
    .a(al_a7b01c14[2]),
    .b(al_85a2bdb0[14]),
    .o(al_f03f7670));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    al_734c4e48 (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_ba3f2ea7),
    .o(al_dfdc4f07));
  AL_MAP_LUT6 #(
    .EQN("(F*~((~B*~(C*~(D*~A))))*~(E)+F*(~B*~(C*~(D*~A)))*~(E)+~(F)*(~B*~(C*~(D*~A)))*E+F*(~B*~(C*~(D*~A)))*E)"),
    .INIT(64'h1303ffff13030000))
    al_410ed209 (
    .a(al_55ed4df1),
    .b(al_f03f7670),
    .c(al_dfdc4f07),
    .d(al_583b2c0d),
    .e(al_8905c135),
    .f(al_25fbce42[46]),
    .o(al_1f3eaa15[14]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_9f7be311 (
    .a(al_f5b7debb),
    .b(al_e2d7fc47),
    .c(al_5fd02584[5]),
    .o(al_8f175a04));
  AL_MAP_LUT6 #(
    .EQN("(~(~(~E*~(~C*~B))*~D)*~(F*~A))"),
    .INIT(64'haa00aaa8ff00fffc))
    al_425290ae (
    .a(al_2ac34e44),
    .b(al_af575898),
    .c(al_bd10bda8),
    .d(al_349edb3b),
    .e(al_792f120f),
    .f(al_4002af45),
    .o(al_dfd548fb));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_61e792d4 (
    .a(al_ba3f2ea7),
    .b(al_f65e6902[7]),
    .o(al_90ba8dd5));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e5561a45 (
    .a(al_653f9409),
    .b(al_7a7cc81),
    .o(al_cee3e376));
  AL_MAP_LUT6 #(
    .EQN("(~F*~(~C*((~B*~A)*~(E)*~(D)+(~B*~A)*E*~(D)+~((~B*~A))*E*D+(~B*~A)*E*D)))"),
    .INIT(64'h00000000f0fefffe))
    al_f2e68434 (
    .a(al_865e8f41),
    .b(al_dfd548fb),
    .c(al_bdf9a7dd),
    .d(al_94dd833a),
    .e(al_90ba8dd5),
    .f(al_cee3e376),
    .o(al_fb22b66));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B))*~(C)+~E*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*~(C)+~(~E)*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*C+~E*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*C)"),
    .INIT(32'h7f4f7040))
    al_1d4c2dd2 (
    .a(al_fb22b66),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[15]),
    .e(al_25fbce42[47]),
    .o(al_1f3eaa15[15]));
  AL_MAP_LUT5 #(
    .EQN("~((~B*A)*~((~E*D))*~(C)+(~B*A)*(~E*D)*~(C)+~((~B*A))*(~E*D)*C+(~B*A)*(~E*D)*C)"),
    .INIT(32'hfdfd0dfd))
    al_c0015280 (
    .a(al_2f34d7b4),
    .b(al_d84a4a58),
    .c(al_e2d7fc47),
    .d(al_5fd02584[7]),
    .e(al_5fd02584[14]),
    .o(al_349edb3b));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    al_8adbb7ff (
    .a(al_ce46ef05),
    .b(al_ba3f2ea7),
    .c(al_3f6865d3),
    .o(al_c6c291a5));
  AL_MAP_LUT6 #(
    .EQN("(A*~(F*~D)*~(E*~C*~B))"),
    .INIT(64'ha800aa00a8a8aaaa))
    al_802493e3 (
    .a(al_c6c291a5),
    .b(al_90d6c009),
    .c(al_c85e3cfa),
    .d(al_65dc271),
    .e(al_8f175a04),
    .f(al_f65e6902[7]),
    .o(al_865e8f41));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(B*(~C*~(E)*~(D)+~C*E*~(D)+~(~C)*E*D+~C*E*D)))"),
    .INIT(32'h11515551))
    al_8bb729ae (
    .a(al_1f0371f8),
    .b(al_7a7cc81),
    .c(al_d84a4a58),
    .d(al_e2d7fc47),
    .e(al_5fd02584[7]),
    .o(al_2ac34e44));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+~(B)*C*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+~(B)*C*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*C*~(D)*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+~(B)*C*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hfcffc0c3f8ffc0c3))
    al_c3052037 (
    .a(al_955e8db5),
    .b(al_843f038d),
    .c(al_ba3f2ea7),
    .d(al_7a7cc81),
    .e(al_47eda15e),
    .f(al_3f6865d3),
    .o(al_f4b0c1c2[16]));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((C*~(B*~A)))*~(D)+~E*(C*~(B*~A))*~(D)+~(~E)*(C*~(B*~A))*D+~E*(C*~(B*~A))*D)"),
    .INIT(32'h4fff4f00))
    al_707fde18 (
    .a(al_9ae3000c),
    .b(al_dec34edc),
    .c(al_5c28a20d),
    .d(al_8905c135),
    .e(al_25fbce42[48]),
    .o(al_1f3eaa15[16]));
  AL_MAP_LUT6 #(
    .EQN("(~E*~((~(A)*~(C)*~(D)*~(F)+A*~(C)*~(D)*~(F)+~(A)*C*~(D)*~(F)+A*C*~(D)*~(F)+~(A)*~(C)*D*~(F)+~(A)*C*~(D)*F+A*C*~(D)*F))*~(B)+~E*(~(A)*~(C)*~(D)*~(F)+A*~(C)*~(D)*~(F)+~(A)*C*~(D)*~(F)+A*C*~(D)*~(F)+~(A)*~(C)*D*~(F)+~(A)*C*~(D)*F+A*C*~(D)*F)*~(B)+~(~E)*(~(A)*~(C)*~(D)*~(F)+A*~(C)*~(D)*~(F)+~(A)*C*~(D)*~(F)+A*C*~(D)*~(F)+~(A)*~(C)*D*~(F)+~(A)*C*~(D)*F+A*C*~(D)*F)*B+~E*(~(A)*~(C)*~(D)*~(F)+A*~(C)*~(D)*~(F)+~(A)*C*~(D)*~(F)+A*C*~(D)*~(F)+~(A)*~(C)*D*~(F)+~(A)*C*~(D)*F+A*C*~(D)*F)*B)"),
    .INIT(64'h00c033f304cc37ff))
    al_73a2e00c (
    .a(al_79632d6f),
    .b(al_ba3f2ea7),
    .c(al_7a7cc81),
    .d(al_47eda15e),
    .e(al_3f6865d3),
    .f(al_55bbd6fb),
    .o(al_5b3d235a));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    al_7072fee8 (
    .a(al_ce46ef05),
    .b(al_c85e3cfa),
    .c(al_4002af45),
    .d(al_47eda15e),
    .o(al_9a488676));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*B)*~C)*~(~D*A))"),
    .INIT(32'hfc54f050))
    al_d95f3d2a (
    .a(al_f4b0c1c2[16]),
    .b(al_5b3d235a),
    .c(al_9a488676),
    .d(al_4002af45),
    .e(al_1f0371f8),
    .o(al_9ae3000c));
  AL_MAP_LUT6 #(
    .EQN("~(E*~((~F*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)))*~(A)+E*(~F*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~(E)*(~F*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*A+E*(~F*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*A)"),
    .INIT(64'haaaaffff028a57df))
    al_7d2387c2 (
    .a(al_a7b01c14[2]),
    .b(al_e2d7fc47),
    .c(al_cf18c1c6[16]),
    .d(al_dc5d601),
    .e(al_85a2bdb0[16]),
    .f(al_653f9409),
    .o(al_5c28a20d));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_2ceecd0 (
    .a(al_4002af45),
    .b(al_843f038d),
    .o(al_94dd833a));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*~(~B*~(~D*~A))))"),
    .INIT(32'h0000f3f2))
    al_b9cff0c7 (
    .a(al_ba6916cf),
    .b(al_357abca7),
    .c(al_d2ba0b0),
    .d(al_4712f186),
    .e(al_bdf9a7dd),
    .o(al_8fddd1ab));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    al_44cd9450 (
    .a(al_653f9409),
    .b(al_e2d7fc47),
    .c(al_cf18c1c6[17]),
    .d(al_39d0a986),
    .o(al_df5cc0b8));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B))*~(D)+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*~(D)+~(~F)*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D)"),
    .INIT(64'hfbffc8fffb00c800))
    al_e0e26cfd (
    .a(al_8fddd1ab),
    .b(al_a7b01c14[2]),
    .c(al_df5cc0b8),
    .d(al_8905c135),
    .e(al_85a2bdb0[17]),
    .f(al_25fbce42[49]),
    .o(al_1f3eaa15[17]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~B*~(~C*~A))"),
    .INIT(32'h00320000))
    al_994c2c9 (
    .a(al_955e8db5),
    .b(al_94dd833a),
    .c(al_792f120f),
    .d(al_ba3f2ea7),
    .e(al_f65e6902[9]),
    .o(al_ba6916cf));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(F*~((E*~(D*A)))*~(C)+F*(E*~(D*A))*~(C)+~(F)*(E*~(D*A))*C+F*(E*~(D*A))*C))"),
    .INIT(64'h2000303023033333))
    al_17add847 (
    .a(al_90d6c009),
    .b(al_ce46ef05),
    .c(al_65dc271),
    .d(al_ba3f2ea7),
    .e(al_3f6865d3),
    .f(al_f65e6902[9]),
    .o(al_357abca7));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    al_22747886 (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_ba3f2ea7),
    .d(al_f65e6902[9]),
    .o(al_d2ba0b0));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D*C)))"),
    .INIT(16'ha888))
    al_8fce3dda (
    .a(al_4002af45),
    .b(al_1f0371f8),
    .c(al_7a7cc81),
    .d(al_f65e6902[9]),
    .o(al_4712f186));
  AL_MAP_LUT5 #(
    .EQN("~((B*~A)*~((E*~D))*~(C)+(B*~A)*(E*~D)*~(C)+~((B*~A))*(E*~D)*C+(B*~A)*(E*~D)*C)"),
    .INIT(32'hfb0bfbfb))
    al_7986ed2a (
    .a(al_e3502e80),
    .b(al_ff37bd99),
    .c(al_e2d7fc47),
    .d(al_5fd02584[12]),
    .e(al_5fd02584[15]),
    .o(al_792f120f));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_65660585 (
    .a(al_a7b01c14[2]),
    .b(al_85a2bdb0[18]),
    .o(al_56afc96e));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)))"),
    .INIT(32'h888aa8aa))
    al_2ece4a24 (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_e2d7fc47),
    .d(al_cf18c1c6[18]),
    .e(al_cf18c1c6[2]),
    .o(al_28a777ae));
  AL_MAP_LUT6 #(
    .EQN("(F*~((~B*~(C*~(~D*~A))))*~(E)+F*(~B*~(C*~(~D*~A)))*~(E)+~(F)*(~B*~(C*~(~D*~A)))*E+F*(~B*~(C*~(~D*~A)))*E)"),
    .INIT(64'h0313ffff03130000))
    al_d3093c79 (
    .a(al_479534eb),
    .b(al_56afc96e),
    .c(al_28a777ae),
    .d(al_bdf9a7dd),
    .e(al_8905c135),
    .f(al_25fbce42[50]),
    .o(al_1f3eaa15[18]));
  AL_MAP_LUT5 #(
    .EQN("(~(C)*~(D)*~((E*~(~B*~A)))+C*~(D)*~((E*~(~B*~A)))+C*D*~((E*~(~B*~A)))+~(C)*~(D)*(E*~(~B*~A))+C*D*(E*~(~B*~A)))"),
    .INIT(32'hf01ff0ff))
    al_72c7c5fd (
    .a(al_955e8db5),
    .b(al_792f120f),
    .c(al_843f038d),
    .d(al_ba3f2ea7),
    .e(al_2d35601b),
    .o(al_77120298));
  AL_MAP_LUT5 #(
    .EQN("(C*B*~(E*~(D*A)))"),
    .INIT(32'h8000c0c0))
    al_2af5b167 (
    .a(al_90d6c009),
    .b(al_65dc271),
    .c(al_1f0371f8),
    .d(al_ba3f2ea7),
    .e(al_3f6865d3),
    .o(al_a32b870b));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*~B))"),
    .INIT(16'h0405))
    al_97cd0e5a (
    .a(al_1f0371f8),
    .b(al_ba3f2ea7),
    .c(al_7a7cc81),
    .d(al_2d35601b),
    .o(al_c96d1fd5));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~((~C*~B))*~(D)+~A*(~C*~B)*~(D)+~(~A)*(~C*~B)*D+~A*(~C*~B)*D)"),
    .INIT(16'hfcaa))
    al_5122bbcb (
    .a(al_77120298),
    .b(al_a32b870b),
    .c(al_c96d1fd5),
    .d(al_4002af45),
    .o(al_479534eb));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_16958d7a (
    .a(al_4002af45),
    .b(al_1f0371f8),
    .o(al_c8e314e6));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((B*A))+D*C*~((B*A))+~(D)*C*(B*A)+D*C*(B*A))"),
    .INIT(16'hf780))
    al_fa7aa239 (
    .a(al_5a744f0f),
    .b(al_6f08d701),
    .c(al_70eedb8b),
    .d(al_85a2bdb0[19]),
    .o(al_d7081cd4));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(~E*C*~(~B*~A)))"),
    .INIT(32'hff00ffe0))
    al_e998760c (
    .a(al_c6dd3893),
    .b(al_b4d3ef2b),
    .c(al_a7b01c14[2]),
    .d(al_d7081cd4),
    .e(al_bdf9a7dd),
    .o(al_704d20e3[19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b1016777 (
    .a(al_704d20e3[19]),
    .b(al_8905c135),
    .c(al_25fbce42[51]),
    .o(al_1f3eaa15[19]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C))"),
    .INIT(16'h08a8))
    al_bd2ac91 (
    .a(al_e22f5efa),
    .b(al_2f34d7b4),
    .c(al_e2d7fc47),
    .d(al_5fd02584[14]),
    .o(al_f2b407ac));
  AL_MAP_LUT6 #(
    .EQN("(C*(B*~(D)*~(E)*~((~F*~A))+~(B)*D*~(E)*~((~F*~A))+B*D*~(E)*~((~F*~A))+~(B)*D*E*~((~F*~A))+B*D*E*~((~F*~A))+B*~(D)*~(E)*(~F*~A)+~(B)*D*~(E)*(~F*~A)+B*D*~(E)*(~F*~A)))"),
    .INIT(64'hf000f0c0a000f0c0))
    al_7aba3eed (
    .a(al_955e8db5),
    .b(al_c8e314e6),
    .c(al_f2b407ac),
    .d(al_e1adfd34),
    .e(al_7a7cc81),
    .f(al_3f6865d3),
    .o(al_c6dd3893));
  AL_MAP_LUT5 #(
    .EQN("(E*B*~(C*~(~D*~A)))"),
    .INIT(32'h0c4c0000))
    al_47fe9e5f (
    .a(al_90d6c009),
    .b(al_1f0371f8),
    .c(al_ba3f2ea7),
    .d(al_7a7cc81),
    .e(al_3f6865d3),
    .o(al_b4d3ef2b));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    al_71d18ce5 (
    .a(al_e2d7fc47),
    .b(al_cf18c1c6[19]),
    .c(al_cf18c1c6[3]),
    .d(al_653f9409),
    .o(al_70eedb8b));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~C*~(~E*~(~D*~B))))"),
    .INIT(32'ha0a0aaa8))
    al_2867ca01 (
    .a(al_a7b01c14[2]),
    .b(al_7c8ae043),
    .c(al_4002af45),
    .d(al_843f038d),
    .e(al_1f0371f8),
    .o(al_2a0680fd));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~A*~(D*~B)))*~(C)+~E*(~A*~(D*~B))*~(C)+~(~E)*(~A*~(D*~B))*C+~E*(~A*~(D*~B))*C)"),
    .INIT(32'hbfafb0a0))
    al_c86cff3b (
    .a(al_2a0680fd),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[1]),
    .e(al_25fbce42[33]),
    .o(al_1f3eaa15[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*~((C*~B)*~((~F*E))*~(D)+(C*~B)*(~F*E)*~(D)+~((C*~B))*(~F*E)*D+(C*~B)*(~F*E)*D))"),
    .INIT(64'haa8aaa8a008aaa8a))
    al_6ba20faa (
    .a(al_78e2749c),
    .b(al_2f34d7b4),
    .c(al_e3502e80),
    .d(al_e2d7fc47),
    .e(al_5fd02584[14]),
    .f(al_5fd02584[15]),
    .o(al_c017beac));
  AL_MAP_LUT6 #(
    .EQN("(F*~C*~A*~(D*~(E*~B)))"),
    .INIT(64'h0105000500000000))
    al_3dcbb3f4 (
    .a(al_96f2b26a),
    .b(al_ac6ff6aa),
    .c(al_d50e9dc4),
    .d(al_4c6b15c2),
    .e(al_57bbe3ad),
    .f(al_653f9409),
    .o(al_f7e849b8));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    al_7d10d813 (
    .a(al_653f9409),
    .b(al_e2d7fc47),
    .c(al_cf18c1c6[20]),
    .d(al_cf18c1c6[4]),
    .o(al_2978bc8a));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B))*~(D)+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*~(D)+~(~F)*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D)"),
    .INIT(64'hfbffc8fffb00c800))
    al_1a77eb6c (
    .a(al_f7e849b8),
    .b(al_a7b01c14[2]),
    .c(al_2978bc8a),
    .d(al_8905c135),
    .e(al_85a2bdb0[20]),
    .f(al_25fbce42[52]),
    .o(al_1f3eaa15[20]));
  AL_MAP_LUT6 #(
    .EQN("(F*~B*~(~E*~D*~C*A))"),
    .INIT(64'h3333333100000000))
    al_45b29bd8 (
    .a(al_75ee8673),
    .b(al_c017beac),
    .c(al_af575898),
    .d(al_7c8ae043),
    .e(al_bd10bda8),
    .f(al_e1adfd34),
    .o(al_96f2b26a));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~D*~(~C*~(E*~A))))"),
    .INIT(32'h33023303))
    al_ce031b9b (
    .a(al_65dc271),
    .b(al_4002af45),
    .c(al_843f038d),
    .d(al_1f0371f8),
    .e(al_78e2749c),
    .o(al_d50e9dc4));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    al_342cf8f2 (
    .a(al_65dc271),
    .b(al_4002af45),
    .c(al_1f0371f8),
    .d(al_78e2749c),
    .o(al_4c6b15c2));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7764f42e (
    .a(al_1f0371f8),
    .b(al_3f6865d3),
    .o(al_57bbe3ad));
  AL_MAP_LUT6 #(
    .EQN("(D*(A*~(B)*~(C)*~(E)*~(F)+~(A)*B*~(C)*~(E)*~(F)+A*B*~(C)*~(E)*~(F)+A*~(B)*C*~(E)*~(F)+~(A)*B*C*~(E)*~(F)+A*B*C*~(E)*~(F)+A*~(B)*~(C)*E*~(F)+A*B*~(C)*E*~(F)+A*~(B)*~(C)*~(E)*F+~(A)*B*~(C)*~(E)*F+A*B*~(C)*~(E)*F+A*~(B)*C*~(E)*F+~(A)*B*C*~(E)*F+A*B*C*~(E)*F+~(A)*~(B)*~(C)*E*F+~(A)*B*~(C)*E*F+~(A)*~(B)*C*E*F+~(A)*B*C*E*F))"),
    .INIT(64'h5500ee000a00ee00))
    al_d234b76b (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_1f0371f8),
    .d(al_f65e6902[3]),
    .e(al_ba3f2ea7),
    .f(al_7a7cc81),
    .o(al_2137298d));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    al_647fe11c (
    .a(al_69efc6c6),
    .b(al_2137298d),
    .c(al_bdf9a7dd),
    .o(al_b0c44f4));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    al_50a02ebe (
    .a(al_653f9409),
    .b(al_e2d7fc47),
    .c(al_cf18c1c6[21]),
    .d(al_cf18c1c6[5]),
    .o(al_da3cc173));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B))*~(D)+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*~(D)+~(~F)*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D)"),
    .INIT(64'hfbffc8fffb00c800))
    al_e0923fba (
    .a(al_b0c44f4),
    .b(al_a7b01c14[2]),
    .c(al_da3cc173),
    .d(al_8905c135),
    .e(al_85a2bdb0[21]),
    .f(al_25fbce42[53]),
    .o(al_1f3eaa15[21]));
  AL_MAP_LUT6 #(
    .EQN("(F*(A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E))"),
    .INIT(64'h55ee4eee00000000))
    al_9cef4712 (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_1f0371f8),
    .d(al_ba3f2ea7),
    .e(al_7a7cc81),
    .f(al_f65e6902[4]),
    .o(al_b931d891));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    al_26d27ad5 (
    .a(al_69efc6c6),
    .b(al_b931d891),
    .c(al_3577d7b9),
    .d(al_55bbd6fb),
    .o(al_1bae5100));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_1b21738f (
    .a(al_a7b01c14[2]),
    .b(al_85a2bdb0[22]),
    .o(al_8bc7d472));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)))"),
    .INIT(32'h888aa8aa))
    al_e6bb6605 (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_e2d7fc47),
    .d(al_cf18c1c6[22]),
    .e(al_cf18c1c6[6]),
    .o(al_55994c98));
  AL_MAP_LUT6 #(
    .EQN("(F*~((~B*~(C*~(~D*~A))))*~(E)+F*(~B*~(C*~(~D*~A)))*~(E)+~(F)*(~B*~(C*~(~D*~A)))*E+F*(~B*~(C*~(~D*~A)))*E)"),
    .INIT(64'h0313ffff03130000))
    al_ffac6b87 (
    .a(al_1bae5100),
    .b(al_8bc7d472),
    .c(al_55994c98),
    .d(al_bdf9a7dd),
    .e(al_8905c135),
    .f(al_25fbce42[54]),
    .o(al_1f3eaa15[22]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_261b85a9 (
    .a(al_90d6c009),
    .b(al_ce46ef05),
    .c(al_c85e3cfa),
    .d(al_3f6865d3),
    .o(al_69efc6c6));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_ed82b986 (
    .a(al_a7b01c14[2]),
    .b(al_85a2bdb0[23]),
    .o(al_136ceed1));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)))"),
    .INIT(32'h888aa8aa))
    al_9b889f83 (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_e2d7fc47),
    .d(al_cf18c1c6[23]),
    .e(al_cf18c1c6[7]),
    .o(al_ffe7e6d4));
  AL_MAP_LUT6 #(
    .EQN("(F*~((~B*~(C*~(~D*~A))))*~(E)+F*(~B*~(C*~(~D*~A)))*~(E)+~(F)*(~B*~(C*~(~D*~A)))*E+F*(~B*~(C*~(~D*~A)))*E)"),
    .INIT(64'h0313ffff03130000))
    al_90a841 (
    .a(al_c51bf9b),
    .b(al_136ceed1),
    .c(al_ffe7e6d4),
    .d(al_bdf9a7dd),
    .e(al_8905c135),
    .f(al_25fbce42[55]),
    .o(al_1f3eaa15[23]));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(~D*~(F*E*C)))"),
    .INIT(64'h8880880088008800))
    al_197a3f08 (
    .a(al_c8e314e6),
    .b(al_65dc271),
    .c(al_7a7cc81),
    .d(al_8f175a04),
    .e(al_2d35601b),
    .f(al_e22f5efa),
    .o(al_a8d5d0d5));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~A*~(~C*~(D*~B))))"),
    .INIT(32'haeaf0000))
    al_12498703 (
    .a(al_843f038d),
    .b(al_1f0371f8),
    .c(al_ba3f2ea7),
    .d(al_7a7cc81),
    .e(al_8f175a04),
    .o(al_4df86c43));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    al_3f354fc1 (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_7a7cc81),
    .d(al_2d35601b),
    .o(al_43099296));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*~A*~(E*D))"),
    .INIT(32'h00010101))
    al_6b6a0df8 (
    .a(al_69efc6c6),
    .b(al_a8d5d0d5),
    .c(al_4df86c43),
    .d(al_43099296),
    .e(al_ba3f2ea7),
    .o(al_c51bf9b));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E*~D*B*~A))"),
    .INIT(32'hf0b0f0f0))
    al_cf374621 (
    .a(al_9e9618ab),
    .b(al_65dc271),
    .c(al_4002af45),
    .d(al_1f0371f8),
    .e(al_55bbd6fb),
    .o(al_343c5862));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B))*~(C)+~E*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*~(C)+~(~E)*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*C+~E*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*C)"),
    .INIT(32'h7f4f7040))
    al_bbd497c0 (
    .a(al_f1e867e0),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[24]),
    .e(al_25fbce42[56]),
    .o(al_1f3eaa15[24]));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~C*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)))"),
    .INIT(32'h30313233))
    al_99e05951 (
    .a(al_90d6c009),
    .b(al_f2b407ac),
    .c(al_c85e3cfa),
    .d(al_3f6865d3),
    .e(al_55bbd6fb),
    .o(al_a683a564));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(E)*~((F*~D))+~(A)*B*~(C)*~(E)*~((F*~D))+A*B*~(C)*~(E)*~((F*~D))+~(A)*~(B)*C*~(E)*~((F*~D))+~(A)*B*C*~(E)*~((F*~D))+A*B*C*~(E)*~((F*~D))+~(A)*~(B)*~(C)*E*~((F*~D))+A*B*~(C)*E*~((F*~D))+~(A)*~(B)*C*E*~((F*~D))+~(A)*B*C*E*~((F*~D))+A*B*C*E*~((F*~D))+~(A)*B*~(C)*~(E)*(F*~D)+A*B*~(C)*~(E)*(F*~D)+~(A)*~(B)*C*~(E)*(F*~D)+~(A)*B*C*~(E)*(F*~D)+A*B*C*~(E)*(F*~D)+A*B*~(C)*E*(F*~D)+~(A)*~(B)*C*E*(F*~D)+~(A)*B*C*E*(F*~D)+A*B*C*E*(F*~D))"),
    .INIT(64'hd9d8dddcd9d9dddd))
    al_d93ae0f0 (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_1f0371f8),
    .d(al_7a7cc81),
    .e(al_55bbd6fb),
    .f(al_e22f5efa),
    .o(al_57675c9b));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_2faf94b7 (
    .a(al_e2d7fc47),
    .b(al_cf18c1c6[24]),
    .c(al_cf18c1c6[8]),
    .o(al_997b23f2));
  AL_MAP_LUT6 #(
    .EQN("(~(~F*~D)*~(~C*~(A*~(E*~B))))"),
    .INIT(64'hf8f8fafaf800fa00))
    al_774f04b0 (
    .a(al_343c5862),
    .b(al_a683a564),
    .c(al_57675c9b),
    .d(al_653f9409),
    .e(al_1f0371f8),
    .f(al_997b23f2),
    .o(al_f1e867e0));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*~(C*~(~E*A))))"),
    .INIT(32'h30331033))
    al_fd09b7af (
    .a(al_f2b407ac),
    .b(al_1f0371f8),
    .c(al_7a7cc81),
    .d(al_3f6865d3),
    .e(al_2d35601b),
    .o(al_a60ca806));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    al_46e1f7b6 (
    .a(al_653f9409),
    .b(al_e2d7fc47),
    .c(al_cf18c1c6[25]),
    .d(al_cf18c1c6[9]),
    .o(al_dffeb202));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~A*~(E*~(C)*~(B)+E*C*~(B)+~(E)*C*B+E*C*B)))*~(D)+~F*(~A*~(E*~(C)*~(B)+E*C*~(B)+~(E)*C*B+E*C*B))*~(D)+~(~F)*(~A*~(E*~(C)*~(B)+E*C*~(B)+~(E)*C*B+E*C*B))*D+~F*(~A*~(E*~(C)*~(B)+E*C*~(B)+~(E)*C*B+E*C*B))*D)"),
    .INIT(64'hfbffeafffb00ea00))
    al_52dd515f (
    .a(al_f57c7577),
    .b(al_a7b01c14[2]),
    .c(al_dffeb202),
    .d(al_8905c135),
    .e(al_85a2bdb0[25]),
    .f(al_25fbce42[57]),
    .o(al_1f3eaa15[25]));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~A*~(~C*~(E)*~(D)+~C*E*~(D)+~(~C)*E*D+~C*E*D)))"),
    .INIT(32'h33232223))
    al_31a9e23f (
    .a(al_843f038d),
    .b(al_ba3f2ea7),
    .c(al_e3502e80),
    .d(al_e2d7fc47),
    .e(al_5fd02584[15]),
    .o(al_370b9296));
  AL_MAP_LUT6 #(
    .EQN("(D*C*~A*~(~E*~(F*~B)))"),
    .INIT(64'h5000100050000000))
    al_a6570b9c (
    .a(al_bdf9a7dd),
    .b(al_370b9296),
    .c(al_5a744f0f),
    .d(al_6f08d701),
    .e(al_4002af45),
    .f(al_3f6865d3),
    .o(al_3cd3cca9));
  AL_MAP_LUT5 #(
    .EQN("~(D*~(C)*~((~(E*B)*~A))+D*C*~((~(E*B)*~A))+~(D)*C*(~(E*B)*~A)+D*C*(~(E*B)*~A))"),
    .INIT(32'h01ef05af))
    al_924833a0 (
    .a(al_c85e3cfa),
    .b(al_47eda15e),
    .c(al_3f6865d3),
    .d(al_78e2749c),
    .e(al_79632d6f),
    .o(al_126b9a65));
  AL_MAP_LUT6 #(
    .EQN("(A*~(D*(B*C*~(E)*~(F)+~(B)*C*E*~(F)+B*C*E*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+B*~(C)*E*F+~(B)*C*E*F+B*C*E*F)))"),
    .INIT(64'h02aa22aa0aaa2aaa))
    al_107f9769 (
    .a(al_3cd3cca9),
    .b(al_a60ca806),
    .c(al_126b9a65),
    .d(al_4002af45),
    .e(al_1f0371f8),
    .f(al_65dc271),
    .o(al_f57c7577));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_bb82e9da (
    .a(al_90d6c009),
    .b(al_c85e3cfa),
    .o(al_73767b69));
  AL_MAP_LUT6 #(
    .EQN("(~B*~((F*~E*~C)*~(A)*~(D)+(F*~E*~C)*A*~(D)+~((F*~E*~C))*A*D+(F*~E*~C)*A*D))"),
    .INIT(64'h1133113011331133))
    al_9f06b678 (
    .a(al_4c1d95c5),
    .b(al_4002af45),
    .c(al_843f038d),
    .d(al_ba3f2ea7),
    .e(al_7a7cc81),
    .f(al_f65e6902[7]),
    .o(al_39ff3661));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((C*~(~D*B*~A)))*~(E)+~F*(C*~(~D*B*~A))*~(E)+~(~F)*(C*~(~D*B*~A))*E+~F*(C*~(~D*B*~A))*E)"),
    .INIT(64'h0f4fffff0f4f0000))
    al_967cac1c (
    .a(al_1c537db1),
    .b(al_dec34edc),
    .c(al_bbb6292e),
    .d(al_39ff3661),
    .e(al_8905c135),
    .f(al_25fbce42[58]),
    .o(al_1f3eaa15[26]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(F*~(C*~(E*~B*A))))"),
    .INIT(64'hd000f000ff00ff00))
    al_239c3347 (
    .a(al_90d6c009),
    .b(al_c85e3cfa),
    .c(al_65dc271),
    .d(al_4002af45),
    .e(al_1f0371f8),
    .f(al_8f175a04),
    .o(al_22e7124d));
  AL_MAP_LUT6 #(
    .EQN("(B*~(~C*~(E*D*~(F*A))))"),
    .INIT(64'hc4c0c0c0ccc0c0c0))
    al_94892913 (
    .a(al_73767b69),
    .b(al_22e7124d),
    .c(al_a60ca806),
    .d(al_349edb3b),
    .e(al_1f0371f8),
    .f(al_3f6865d3),
    .o(al_1c537db1));
  AL_MAP_LUT6 #(
    .EQN("~(F*~((~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)))*~(A)+F*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*~(A)+~(F)*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A+F*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A)"),
    .INIT(64'h888aa8aadddffdff))
    al_8ba6922e (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_e2d7fc47),
    .d(al_cf18c1c6[26]),
    .e(al_cf18c1c6[10]),
    .f(al_85a2bdb0[26]),
    .o(al_bbb6292e));
  AL_MAP_LUT5 #(
    .EQN("(C*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(A)+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)+~(C)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A)"),
    .INIT(32'hfad87250))
    al_1435a3 (
    .a(al_843f038d),
    .b(al_7a7cc81),
    .c(al_8f175a04),
    .d(al_78e2749c),
    .e(al_f65e6902[7]),
    .o(al_4c1d95c5));
  AL_MAP_LUT6 #(
    .EQN("(C*~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(F)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*F*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*F*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*F*B))"),
    .INIT(64'h00201030c0e0d0f0))
    al_60339c44 (
    .a(al_90d6c009),
    .b(al_c85e3cfa),
    .c(al_1f0371f8),
    .d(al_f65e6902[3]),
    .e(al_3f6865d3),
    .f(al_55bbd6fb),
    .o(al_ea06ea2d));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5f7aff7f))
    al_68774070 (
    .a(al_843f038d),
    .b(al_f65e6902[3]),
    .c(al_ba3f2ea7),
    .d(al_7a7cc81),
    .e(al_47eda15e),
    .o(al_8b49a361));
  AL_MAP_LUT6 #(
    .EQN("~(~C*~((~A*~(B*~(F*~D))))*~(E)+~C*(~A*~(B*~(F*~D)))*~(E)+~(~C)*(~A*~(B*~(F*~D)))*E+~C*(~A*~(B*~(F*~D)))*E)"),
    .INIT(64'heeaaf0f0eeeef0f0))
    al_73551ffa (
    .a(al_ea06ea2d),
    .b(al_a60ca806),
    .c(al_8b49a361),
    .d(al_65dc271),
    .e(al_4002af45),
    .f(al_55bbd6fb),
    .o(al_dccb8299));
  AL_MAP_LUT6 #(
    .EQN("~(F*~((~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)))*~(A)+F*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*~(A)+~(F)*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A+F*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A)"),
    .INIT(64'h888aa8aadddffdff))
    al_16c9549c (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_e2d7fc47),
    .d(al_cf18c1c6[27]),
    .e(al_cf18c1c6[11]),
    .f(al_85a2bdb0[27]),
    .o(al_bd675004));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((C*~(B*~A)))*~(D)+~E*(C*~(B*~A))*~(D)+~(~E)*(C*~(B*~A))*D+~E*(C*~(B*~A))*D)"),
    .INIT(32'h4fff4f00))
    al_f6c8fd5b (
    .a(al_dccb8299),
    .b(al_dec34edc),
    .c(al_bd675004),
    .d(al_8905c135),
    .e(al_25fbce42[59]),
    .o(al_1f3eaa15[27]));
  AL_MAP_LUT6 #(
    .EQN("(B*(A*~((E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D))*~(C)+A*(E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)*~(C)+~(A)*(E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)*C+A*(E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)*C))"),
    .INIT(64'hc8c8c80808c80808))
    al_da98dd8e (
    .a(al_7aa9f4ee[31]),
    .b(al_4002af45),
    .c(al_843f038d),
    .d(al_e2d7fc47),
    .e(al_cf18c1c6[31]),
    .f(al_cf18c1c6[15]),
    .o(al_8778492e[31]));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D)*~((~B*A))+C*D*~((~B*A))+~(C)*D*(~B*A)+C*D*(~B*A))"),
    .INIT(16'h0d2f))
    al_2d86f2c8 (
    .a(al_90d6c009),
    .b(al_7a7cc81),
    .c(al_3f6865d3),
    .d(al_f65e6902[4]),
    .o(al_3e7bf97e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hca00cacffa30faff))
    al_7e0326d6 (
    .a(al_3e7bf97e),
    .b(al_3577d7b9),
    .c(al_ce46ef05),
    .d(al_ba3f2ea7),
    .e(al_f65e6902[9]),
    .f(al_8778492e[31]),
    .o(al_e99a5572));
  AL_MAP_LUT6 #(
    .EQN("~(F*~((~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)))*~(A)+F*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*~(A)+~(F)*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A+F*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A)"),
    .INIT(64'h888aa8aadddffdff))
    al_2bf77470 (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_e2d7fc47),
    .d(al_cf18c1c6[28]),
    .e(al_cf18c1c6[12]),
    .f(al_85a2bdb0[28]),
    .o(al_47e27082));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((C*~(B*~A)))*~(D)+~E*(C*~(B*~A))*~(D)+~(~E)*(C*~(B*~A))*D+~E*(C*~(B*~A))*D)"),
    .INIT(32'h4fff4f00))
    al_d4da34c3 (
    .a(al_e99a5572),
    .b(al_dec34edc),
    .c(al_47e27082),
    .d(al_8905c135),
    .e(al_25fbce42[60]),
    .o(al_1f3eaa15[28]));
  AL_MAP_LUT6 #(
    .EQN("~(F*~((~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)))*~(A)+F*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*~(A)+~(F)*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A+F*(~B*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A)"),
    .INIT(64'h888aa8aadddffdff))
    al_c29ece0c (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_e2d7fc47),
    .d(al_cf18c1c6[29]),
    .e(al_cf18c1c6[13]),
    .f(al_85a2bdb0[29]),
    .o(al_b9001309));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h5f5f03135f5fff5f))
    al_bc48cc9 (
    .a(al_7aa9f4ee[31]),
    .b(al_3577d7b9),
    .c(al_4002af45),
    .d(al_1f0371f8),
    .e(al_ba3f2ea7),
    .f(al_2d35601b),
    .o(al_d56de4dc));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((B*~(~C*A)))*~(D)+~E*(B*~(~C*A))*~(D)+~(~E)*(B*~(~C*A))*D+~E*(B*~(~C*A))*D)"),
    .INIT(32'h3bff3b00))
    al_a1c396a8 (
    .a(al_dec34edc),
    .b(al_b9001309),
    .c(al_d56de4dc),
    .d(al_8905c135),
    .e(al_25fbce42[61]),
    .o(al_1f3eaa15[29]));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*((D*C)*~(F)*~(E)+(D*C)*F*~(E)+~((D*C))*F*E+(D*C)*F*E))"),
    .INIT(64'h4444400000004000))
    al_71b537bf (
    .a(al_4aed8be6),
    .b(al_47eda15e),
    .c(al_d84a4a58),
    .d(al_c524b83f),
    .e(al_e2d7fc47),
    .f(al_88242571),
    .o(al_90d6c009));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    al_1d597cf7 (
    .a(al_90d6c009),
    .b(al_ba3f2ea7),
    .c(al_7a7cc81),
    .o(al_ac6ff6aa));
  AL_MAP_LUT6 #(
    .EQN("(~C*~(~(F*~D*B)*~(~E*~A)))"),
    .INIT(64'h000c050d00000505))
    al_1af2545f (
    .a(al_ac6ff6aa),
    .b(al_695857c1),
    .c(al_bdf9a7dd),
    .d(al_75ee8673),
    .e(al_ce46ef05),
    .f(al_e1adfd34),
    .o(al_31e9afe8));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_56eac5ab (
    .a(al_653f9409),
    .b(al_78e2749c),
    .o(al_575fad37));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B))*~(D)+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*~(D)+~(~F)*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D)"),
    .INIT(64'hfbffc8fffb00c800))
    al_98ceb2fd (
    .a(al_31e9afe8),
    .b(al_a7b01c14[2]),
    .c(al_575fad37),
    .d(al_8905c135),
    .e(al_85a2bdb0[2]),
    .f(al_25fbce42[34]),
    .o(al_1f3eaa15[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_5e3e5055 (
    .a(al_5fd02584[0]),
    .b(al_5fd02584[13]),
    .o(al_ec9911d2));
  AL_MAP_LUT6 #(
    .EQN("~((~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*~(F)*~(C)+(~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*F*~(C)+~((~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)))*F*C+(~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*F*C)"),
    .INIT(64'h0c0e0d0ffcfefdff))
    al_30ab7da4 (
    .a(al_a0b8db17),
    .b(al_c6ff495c),
    .c(al_e2d7fc47),
    .d(al_cf18c1c6[29]),
    .e(al_cf18c1c6[13]),
    .f(al_ec9911d2),
    .o(al_ce46ef05));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_a82d2a37 (
    .a(al_a8af8112),
    .b(al_e2d7fc47),
    .c(al_5fd02584[2]),
    .o(al_78e2749c));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_e2f4c44f (
    .a(al_77bf7190),
    .b(al_e2d7fc47),
    .c(al_5fd02584[1]),
    .o(al_e1adfd34));
  AL_MAP_LUT6 #(
    .EQN("(D*~(C*~B*~A*~(F*~E)))"),
    .INIT(64'hef00ff00ef00ef00))
    al_346d4be3 (
    .a(al_1f0371f8),
    .b(al_ba3f2ea7),
    .c(al_7a7cc81),
    .d(al_3f6865d3),
    .e(al_2d35601b),
    .f(al_e22f5efa),
    .o(al_7aa9f4ee[31]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_bdc2e628 (
    .a(al_4002af45),
    .b(al_843f038d),
    .o(al_583b2c0d));
  AL_MAP_LUT5 #(
    .EQN("(D*C*A*~(E*B))"),
    .INIT(32'h2000a000))
    al_7ed537d7 (
    .a(al_c7467d2d),
    .b(al_bd10bda8),
    .c(al_7a7cc81),
    .d(al_2d35601b),
    .e(al_e22f5efa),
    .o(al_abfe390c));
  AL_MAP_LUT6 #(
    .EQN("(C*~(~A*~(B*~(F)*~((~E*D))+B*F*~((~E*D))+~(B)*F*(~E*D)+B*F*(~E*D))))"),
    .INIT(64'he0e0f0e0e0e0a0e0))
    al_6f104752 (
    .a(al_abfe390c),
    .b(al_7aa9f4ee[31]),
    .c(al_583b2c0d),
    .d(al_1f0371f8),
    .e(al_ba3f2ea7),
    .f(al_47eda15e),
    .o(al_da123ab6));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    al_a772da51 (
    .a(al_653f9409),
    .b(al_e2d7fc47),
    .c(al_cf18c1c6[30]),
    .d(al_cf18c1c6[14]),
    .o(al_f92423e));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B))*~(D)+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*~(D)+~(~F)*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D)"),
    .INIT(64'hfbffc8fffb00c800))
    al_634b7cac (
    .a(al_da123ab6),
    .b(al_a7b01c14[2]),
    .c(al_f92423e),
    .d(al_8905c135),
    .e(al_85a2bdb0[30]),
    .f(al_25fbce42[62]),
    .o(al_1f3eaa15[30]));
  AL_MAP_LUT5 #(
    .EQN("(E*~((D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))*~(C)+E*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*~(C)+~(E)*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C+E*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C)"),
    .INIT(32'hbf8fb080))
    al_589f1b34 (
    .a(al_8778492e[31]),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[31]),
    .e(al_25fbce42[63]),
    .o(al_1f3eaa15[31]));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((~D*~B))*~(A)+C*(~D*~B)*~(A)+~(C)*(~D*~B)*A+C*(~D*~B)*A)"),
    .INIT(16'haf8d))
    al_f11a5e9a (
    .a(al_653f9409),
    .b(al_ce46ef05),
    .c(al_f65e6902[3]),
    .d(al_ba3f2ea7),
    .o(al_b4ed90bc));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B))*~(C)+~E*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*~(C)+~(~E)*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*C+~E*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B)*C)"),
    .INIT(32'h7f4f7040))
    al_9ec74988 (
    .a(al_b4ed90bc),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[3]),
    .e(al_25fbce42[35]),
    .o(al_1f3eaa15[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_63c61a3c (
    .a(iBusAhb_HRDATA[23]),
    .b(al_b86dd14b[24]),
    .c(al_d518b626),
    .o(al_cf18c1c6[23]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_ef6d881c (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[28]),
    .c(al_cf18c1c6[12]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_ff37bd99));
  AL_MAP_LUT5 #(
    .EQN("~((~B*A)*~((E*~D))*~(C)+(~B*A)*(E*~D)*~(C)+~((~B*A))*(E*~D)*C+(~B*A)*(E*~D)*C)"),
    .INIT(32'hfd0dfdfd))
    al_7652d595 (
    .a(al_97cb05f),
    .b(al_ff37bd99),
    .c(al_e2d7fc47),
    .d(al_5fd02584[8]),
    .e(al_5fd02584[12]),
    .o(al_b0110a42));
  AL_MAP_LUT6 #(
    .EQN("(~B*~A*((D*C)*~(F)*~(E)+(D*C)*F*~(E)+~((D*C))*F*E+(D*C)*F*E))"),
    .INIT(64'h1111100000001000))
    al_7f5da429 (
    .a(al_4aed8be6),
    .b(al_b0110a42),
    .c(al_d84a4a58),
    .d(al_c524b83f),
    .e(al_e2d7fc47),
    .f(al_88242571),
    .o(al_75ee8673));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*~(~C*~B*~A)))"),
    .INIT(32'h01ff0000))
    al_52982dd1 (
    .a(al_75ee8673),
    .b(al_af575898),
    .c(al_bd10bda8),
    .d(al_843f038d),
    .e(al_7a7cc81),
    .o(al_33012db3));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff44cf440044cf44))
    al_aa256713 (
    .a(al_33012db3),
    .b(al_c7467d2d),
    .c(al_c85e3cfa),
    .d(al_4002af45),
    .e(al_843f038d),
    .f(al_f65e6902[4]),
    .o(al_8778492e[4]));
  AL_MAP_LUT5 #(
    .EQN("(E*~((D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))*~(C)+E*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*~(C)+~(E)*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C+E*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C)"),
    .INIT(32'hbf8fb080))
    al_7f61344f (
    .a(al_8778492e[4]),
    .b(al_a7b01c14[2]),
    .c(al_8905c135),
    .d(al_85a2bdb0[4]),
    .e(al_25fbce42[36]),
    .o(al_1f3eaa15[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ca71f874 (
    .a(iBusAhb_HRDATA[28]),
    .b(al_b86dd14b[29]),
    .c(al_d518b626),
    .o(al_cf18c1c6[28]));
  AL_MAP_LUT5 #(
    .EQN("~((B*A)*~((~E*~D))*~(C)+(B*A)*(~E*~D)*~(C)+~((B*A))*(~E*~D)*C+(B*A)*(~E*~D)*C)"),
    .INIT(32'hf7f7f707))
    al_e8f3294b (
    .a(al_d344e0e5),
    .b(al_87b30ed5),
    .c(al_e2d7fc47),
    .d(al_5fd02584[10]),
    .e(al_5fd02584[11]),
    .o(al_4aed8be6));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7aecd360 (
    .a(iBusAhb_HRDATA[7]),
    .b(al_b86dd14b[8]),
    .c(al_d518b626),
    .o(al_cf18c1c6[7]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_8c170a3a (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[23]),
    .c(al_cf18c1c6[7]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_d84a4a58));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_8d9a670 (
    .a(al_5fd02584[7]),
    .b(al_5fd02584[9]),
    .o(al_88242571));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_817d98c6 (
    .a(iBusAhb_HRDATA[12]),
    .b(al_b86dd14b[13]),
    .c(al_d518b626),
    .o(al_cf18c1c6[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_4b71ebdf (
    .a(al_7a7cc81),
    .b(al_2d35601b),
    .c(al_e22f5efa),
    .o(al_9e9618ab));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((~D*~A))*~(E)*~(F)+~(B)*C*~((~D*~A))*~(E)*~(F)+~(B)*~(C)*(~D*~A)*~(E)*~(F)+B*~(C)*(~D*~A)*~(E)*~(F)+~(B)*C*(~D*~A)*~(E)*~(F)+B*C*(~D*~A)*~(E)*~(F)+~(B)*~(C)*~((~D*~A))*E*~(F)+~(B)*C*~((~D*~A))*E*~(F)+~(B)*~(C)*(~D*~A)*E*~(F)+B*~(C)*(~D*~A)*E*~(F)+~(B)*C*(~D*~A)*E*~(F)+B*C*(~D*~A)*E*~(F)+~(B)*~(C)*~((~D*~A))*~(E)*F+~(B)*~(C)*(~D*~A)*~(E)*F+B*~(C)*(~D*~A)*~(E)*F+B*C*(~D*~A)*~(E)*F)"),
    .INIT(64'h0000034733773377))
    al_d35e2dce (
    .a(al_9e9618ab),
    .b(al_4002af45),
    .c(al_843f038d),
    .d(al_1f0371f8),
    .e(al_ba3f2ea7),
    .f(al_7a7cc81),
    .o(al_c74661));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*~A*~(~E*D))"),
    .INIT(32'h04040004))
    al_8bb9eebf (
    .a(al_c74661),
    .b(al_a7b01c14[2]),
    .c(al_bdf9a7dd),
    .d(al_90d6c009),
    .e(al_c85e3cfa),
    .o(al_387eb97));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h8adf))
    al_a68ba363 (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_8f175a04),
    .d(al_85a2bdb0[5]),
    .o(al_d7a80970));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*~A))*~(C)+~D*(B*~A)*~(C)+~(~D)*(B*~A)*C+~D*(B*~A)*C)"),
    .INIT(16'hbfb0))
    al_1b2461ef (
    .a(al_387eb97),
    .b(al_d7a80970),
    .c(al_8905c135),
    .d(al_25fbce42[37]),
    .o(al_1f3eaa15[5]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*B*A)"),
    .INIT(32'h08000000))
    al_5bf48d76 (
    .a(al_955e8db5),
    .b(al_c7467d2d),
    .c(al_4002af45),
    .d(al_843f038d),
    .e(al_7a7cc81),
    .o(al_14c6d47a));
  AL_MAP_LUT5 #(
    .EQN("(C*((B*~A)*~(E)*~(D)+(B*~A)*E*~(D)+~((B*~A))*E*D+(B*~A)*E*D))"),
    .INIT(32'hf0400040))
    al_46ba149e (
    .a(al_c7467d2d),
    .b(al_c85e3cfa),
    .c(al_4002af45),
    .d(al_843f038d),
    .e(al_55bbd6fb),
    .o(al_d63f10c0));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*~((~B*~A))*~(C)+~E*(~B*~A)*~(C)+~(~E)*(~B*~A)*C+~E*(~B*~A)*C))*~(D)+~F*(~E*~((~B*~A))*~(C)+~E*(~B*~A)*~(C)+~(~E)*(~B*~A)*C+~E*(~B*~A)*C)*~(D)+~(~F)*(~E*~((~B*~A))*~(C)+~E*(~B*~A)*~(C)+~(~E)*(~B*~A)*C+~E*(~B*~A)*C)*D+~F*(~E*~((~B*~A))*~(C)+~E*(~B*~A)*~(C)+~(~E)*(~B*~A)*C+~E*(~B*~A)*C)*D)"),
    .INIT(64'hefffe0ffef00e000))
    al_70fac76 (
    .a(al_14c6d47a),
    .b(al_d63f10c0),
    .c(al_a7b01c14[2]),
    .d(al_8905c135),
    .e(al_85a2bdb0[6]),
    .f(al_25fbce42[38]),
    .o(al_1f3eaa15[6]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_2ba8f856 (
    .a(al_ff37bd99),
    .b(al_e2d7fc47),
    .c(al_5fd02584[12]),
    .o(al_3f6865d3));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    al_e13c5581 (
    .a(al_79632d6f),
    .b(al_47eda15e),
    .c(al_3f6865d3),
    .o(al_12790a23));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf400f7ff))
    al_fa9d2cb (
    .a(al_12790a23),
    .b(al_955e8db5),
    .c(al_ba3f2ea7),
    .d(al_7a7cc81),
    .e(al_f65e6902[7]),
    .o(al_c115942c));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E*~((C*~B))*~(A)+E*(C*~B)*~(A)+~(E)*(C*~B)*A+E*(C*~B)*A))"),
    .INIT(32'h8a00df00))
    al_b168891 (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_f65e6902[7]),
    .d(al_8905c135),
    .e(al_85a2bdb0[7]),
    .o(al_d68a240f));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*C*D*E)"),
    .INIT(32'h20e03dfd))
    al_e4360128 (
    .a(al_1f0371f8),
    .b(al_ba3f2ea7),
    .c(al_7a7cc81),
    .d(al_3f6865d3),
    .e(al_f65e6902[7]),
    .o(al_3ce9d83));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    al_93a89af8 (
    .a(al_3ce9d83),
    .b(al_3577d7b9),
    .c(al_4002af45),
    .d(al_78e2749c),
    .o(al_19463fbe));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_c2b6c3fd (
    .a(al_8905c135),
    .b(al_25fbce42[39]),
    .o(al_ef0a8112));
  AL_MAP_LUT6 #(
    .EQN("(~F*~(C*~(B*~(D*~(E*~A)))))"),
    .INIT(64'h000000004fcf0fcf))
    al_6059ce6f (
    .a(al_c115942c),
    .b(al_dec34edc),
    .c(al_d68a240f),
    .d(al_19463fbe),
    .e(al_e1adfd34),
    .f(al_ef0a8112),
    .o(al_1f3eaa15[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_7245d745 (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_7a7cc81),
    .o(al_3577d7b9));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5cdb973a (
    .a(al_a7b01c14[2]),
    .b(al_bdf9a7dd),
    .o(al_dec34edc));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_83f813ca (
    .a(al_d84a4a58),
    .b(al_e2d7fc47),
    .c(al_5fd02584[7]),
    .o(al_f65e6902[7]));
  AL_MAP_LUT5 #(
    .EQN("(~A*((C*B)*~(E)*~(D)+(C*B)*E*~(D)+~((C*B))*E*D+(C*B)*E*D))"),
    .INIT(32'h55400040))
    al_763f9554 (
    .a(al_4aed8be6),
    .b(al_d84a4a58),
    .c(al_c524b83f),
    .d(al_e2d7fc47),
    .e(al_88242571),
    .o(al_79632d6f));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_813a0f4a (
    .a(iBusAhb_HRDATA[31]),
    .b(al_b86dd14b[32]),
    .c(al_d518b626),
    .o(al_cf18c1c6[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9980b71b (
    .a(al_f56de171),
    .b(al_bccf82af),
    .c(al_bd9d7d67),
    .o(al_e2d7fc47));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~((~D*~C))*~(A)+~B*(~D*~C)*~(A)+~(~B)*(~D*~C)*A+~B*(~D*~C)*A)"),
    .INIT(16'heee4))
    al_ed0f5519 (
    .a(al_bd9d7d67),
    .b(al_a2250ee),
    .c(al_9c16c2f5),
    .d(al_126b3afd[1]),
    .o(al_a0b8db17));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d1d5a59d (
    .a(iBusAhb_HRDATA[8]),
    .b(al_b86dd14b[9]),
    .c(al_d518b626),
    .o(al_cf18c1c6[8]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_c0e15a6 (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[24]),
    .c(al_cf18c1c6[8]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_97cb05f));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_dc82c151 (
    .a(al_97cb05f),
    .b(al_e2d7fc47),
    .c(al_5fd02584[8]),
    .o(al_47eda15e));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_4c07502f (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[16]),
    .c(al_dc5d601),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_c6ff495c));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9472ccc1 (
    .a(iBusAhb_HRDATA[13]),
    .b(al_b86dd14b[14]),
    .c(al_d518b626),
    .o(al_cf18c1c6[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9f9a1d4 (
    .a(iBusAhb_HRDATA[30]),
    .b(al_b86dd14b[31]),
    .c(al_d518b626),
    .o(al_cf18c1c6[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_230d7614 (
    .a(iBusAhb_HRDATA[14]),
    .b(al_b86dd14b[15]),
    .c(al_d518b626),
    .o(al_cf18c1c6[14]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_f249aeb (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[30]),
    .c(al_cf18c1c6[14]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_2f34d7b4));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8046ac9 (
    .a(iBusAhb_HRDATA[15]),
    .b(al_b86dd14b[16]),
    .c(al_d518b626),
    .o(al_cf18c1c6[15]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_97d91b30 (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[31]),
    .c(al_cf18c1c6[15]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_e3502e80));
  AL_MAP_LUT5 #(
    .EQN("~((B*~A)*~((~E*D))*~(C)+(B*~A)*(~E*D)*~(C)+~((B*~A))*(~E*D)*C+(B*~A)*(~E*D)*C)"),
    .INIT(32'hfbfb0bfb))
    al_50799445 (
    .a(al_2f34d7b4),
    .b(al_e3502e80),
    .c(al_e2d7fc47),
    .d(al_5fd02584[14]),
    .e(al_5fd02584[15]),
    .o(al_c85e3cfa));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_122ec21b (
    .a(al_c6ff495c),
    .b(al_e2d7fc47),
    .c(al_5fd02584[0]),
    .o(al_4002af45));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_7e48c805 (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[17]),
    .c(al_39d0a986),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_77bf7190));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_249f92fc (
    .a(iBusAhb_HRDATA[18]),
    .b(al_b86dd14b[19]),
    .c(al_d518b626),
    .o(al_cf18c1c6[18]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_27808921 (
    .a(al_77bf7190),
    .b(al_e2d7fc47),
    .c(al_5fd02584[1]),
    .o(al_843f038d));
  AL_MAP_LUT5 #(
    .EQN("((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*~(E)*~(B)+(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*E*~(B)+~((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))*E*B+(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*E*B)"),
    .INIT(32'hfdec3120))
    al_b5c4a146 (
    .a(al_a0b8db17),
    .b(al_e2d7fc47),
    .c(al_cf18c1c6[29]),
    .d(al_cf18c1c6[13]),
    .e(al_5fd02584[13]),
    .o(al_1f0371f8));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d94944fe (
    .a(iBusAhb_HRDATA[3]),
    .b(al_b86dd14b[4]),
    .c(al_d518b626),
    .o(al_cf18c1c6[3]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_7feb057c (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[19]),
    .c(al_cf18c1c6[3]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_31f2e639));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_1c958593 (
    .a(al_31f2e639),
    .b(al_e2d7fc47),
    .c(al_5fd02584[3]),
    .o(al_f65e6902[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_1daf24b7 (
    .a(al_2f34d7b4),
    .b(al_e2d7fc47),
    .c(al_5fd02584[14]),
    .o(al_ba3f2ea7));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a8ac762d (
    .a(iBusAhb_HRDATA[19]),
    .b(al_b86dd14b[20]),
    .c(al_d518b626),
    .o(al_cf18c1c6[19]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_4af5ee88 (
    .a(al_e3502e80),
    .b(al_e2d7fc47),
    .c(al_5fd02584[15]),
    .o(al_7a7cc81));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4d9bf963 (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_1f0371f8),
    .o(al_bdf9a7dd));
  AL_MAP_LUT5 #(
    .EQN("~((~B*~A)*~((E*D))*~(C)+(~B*~A)*(E*D)*~(C)+~((~B*~A))*(E*D)*C+(~B*~A)*(E*D)*C)"),
    .INIT(32'h0efefefe))
    al_f756fbe6 (
    .a(al_c6ff495c),
    .b(al_77bf7190),
    .c(al_e2d7fc47),
    .d(al_5fd02584[0]),
    .e(al_5fd02584[1]),
    .o(al_653f9409));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8ad08eed (
    .a(iBusAhb_HRDATA[5]),
    .b(al_b86dd14b[6]),
    .c(al_d518b626),
    .o(al_cf18c1c6[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5ceb8ebc (
    .a(iBusAhb_HRDATA[4]),
    .b(al_b86dd14b[5]),
    .c(al_d518b626),
    .o(al_cf18c1c6[4]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_9a4f67dd (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[20]),
    .c(al_cf18c1c6[4]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_3629238d));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ee0ced7 (
    .a(iBusAhb_HRDATA[20]),
    .b(al_b86dd14b[21]),
    .c(al_d518b626),
    .o(al_cf18c1c6[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_500e185e (
    .a(iBusAhb_HRDATA[6]),
    .b(al_b86dd14b[7]),
    .c(al_d518b626),
    .o(al_cf18c1c6[6]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_bec83b0a (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[22]),
    .c(al_cf18c1c6[6]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_12584de1));
  AL_MAP_LUT5 #(
    .EQN("~((~B*~A)*~((E*D))*~(C)+(~B*~A)*(E*D)*~(C)+~((~B*~A))*(E*D)*C+(~B*~A)*(E*D)*C)"),
    .INIT(32'h0efefefe))
    al_2717b04a (
    .a(al_2f34d7b4),
    .b(al_e3502e80),
    .c(al_e2d7fc47),
    .d(al_5fd02584[14]),
    .e(al_5fd02584[15]),
    .o(al_65dc271));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_58b527a8 (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[21]),
    .c(al_cf18c1c6[5]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_f5b7debb));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_c4b4ed56 (
    .a(al_5c72a609[0]),
    .b(al_5c72a609[1]),
    .c(al_5c72a609[2]),
    .o(al_8905c135));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1063e022 (
    .a(iBusAhb_HRDATA[2]),
    .b(al_b86dd14b[3]),
    .c(al_d518b626),
    .o(al_cf18c1c6[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3b335986 (
    .a(iBusAhb_HRDATA[21]),
    .b(al_b86dd14b[22]),
    .c(al_d518b626),
    .o(al_cf18c1c6[21]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_1aace9ed (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[18]),
    .c(al_cf18c1c6[2]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_a8af8112));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_6a20d836 (
    .a(al_5fd02584[2]),
    .b(al_5fd02584[3]),
    .c(al_5fd02584[4]),
    .o(al_42488c02));
  AL_MAP_LUT5 #(
    .EQN("~((C*B*A)*~(E)*~(D)+(C*B*A)*E*~(D)+~((C*B*A))*E*D+(C*B*A)*E*D)"),
    .INIT(32'h007fff7f))
    al_54db4c1a (
    .a(al_31f2e639),
    .b(al_3629238d),
    .c(al_a8af8112),
    .d(al_e2d7fc47),
    .e(al_42488c02),
    .o(al_af575898));
  AL_MAP_LUT5 #(
    .EQN("~((B*A)*~((~E*~D))*~(C)+(B*A)*(~E*~D)*~(C)+~((B*A))*(~E*~D)*C+(B*A)*(~E*~D)*C)"),
    .INIT(32'hf7f7f707))
    al_860e1f0e (
    .a(al_12584de1),
    .b(al_f5b7debb),
    .c(al_e2d7fc47),
    .d(al_5fd02584[5]),
    .e(al_5fd02584[6]),
    .o(al_bd10bda8));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_e4cd358b (
    .a(al_af575898),
    .b(al_bd10bda8),
    .o(al_955e8db5));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_15265a22 (
    .a(al_1f0371f8),
    .b(al_ba3f2ea7),
    .o(al_c7467d2d));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b456eaf1 (
    .a(iBusAhb_HRDATA[22]),
    .b(al_b86dd14b[23]),
    .c(al_d518b626),
    .o(al_cf18c1c6[22]));
  AL_MAP_LUT5 #(
    .EQN("(E*C*B*~(D*A))"),
    .INIT(32'h40c00000))
    al_4d09ab69 (
    .a(al_955e8db5),
    .b(al_65dc271),
    .c(al_843f038d),
    .d(al_7a7cc81),
    .e(al_47eda15e),
    .o(al_e240543c));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E*~C)*~(F*~(B*~A)))"),
    .INIT(64'h40004400f000ff00))
    al_ef1b7545 (
    .a(al_c7467d2d),
    .b(al_c85e3cfa),
    .c(al_65dc271),
    .d(al_4002af45),
    .e(al_f65e6902[3]),
    .f(al_47eda15e),
    .o(al_88a18e08));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*~B))"),
    .INIT(16'h5545))
    al_afb9d7a (
    .a(al_4002af45),
    .b(al_843f038d),
    .c(al_f65e6902[3]),
    .d(al_7a7cc81),
    .o(al_1754eacf));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*~A))"),
    .INIT(16'h0023))
    al_75aaa46b (
    .a(al_e240543c),
    .b(al_88a18e08),
    .c(al_1754eacf),
    .d(al_bdf9a7dd),
    .o(al_a72e375d));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b6e71ff8 (
    .a(al_653f9409),
    .b(al_47eda15e),
    .o(al_2df3af97));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_15bdf64a (
    .a(iBusAhb_HRDATA[24]),
    .b(al_b86dd14b[25]),
    .c(al_d518b626),
    .o(al_cf18c1c6[24]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B))*~(D)+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*~(D)+~(~F)*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D+~F*(~E*~((~C*~A))*~(B)+~E*(~C*~A)*~(B)+~(~E)*(~C*~A)*B+~E*(~C*~A)*B)*D)"),
    .INIT(64'hfbffc8fffb00c800))
    al_db6104d5 (
    .a(al_a72e375d),
    .b(al_a7b01c14[2]),
    .c(al_2df3af97),
    .d(al_8905c135),
    .e(al_85a2bdb0[8]),
    .f(al_25fbce42[40]),
    .o(al_1f3eaa15[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_505eaf59 (
    .a(iBusAhb_HRDATA[29]),
    .b(al_b86dd14b[30]),
    .c(al_d518b626),
    .o(al_cf18c1c6[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_29c8455e (
    .a(iBusAhb_HRDATA[25]),
    .b(al_b86dd14b[26]),
    .c(al_d518b626),
    .o(al_cf18c1c6[25]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_993ef97f (
    .a(al_c524b83f),
    .b(al_e2d7fc47),
    .c(al_5fd02584[9]),
    .o(al_f65e6902[9]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_d8e6e91f (
    .a(al_af575898),
    .b(al_7c8ae043),
    .c(al_bd10bda8),
    .o(al_695857c1));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    al_b9927015 (
    .a(al_a7b01c14[2]),
    .b(al_653f9409),
    .c(al_f65e6902[9]),
    .o(al_7244a2ec));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    al_31bfbe99 (
    .a(al_a7b01c14[2]),
    .b(al_8905c135),
    .c(al_85a2bdb0[9]),
    .o(al_52be31ea));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*A))*~(B)+C*(D*A)*~(B)+~(C)*(D*A)*B+C*(D*A)*B)"),
    .INIT(16'h47cf))
    al_1f7c0981 (
    .a(al_ba3f2ea7),
    .b(al_7a7cc81),
    .c(al_f65e6902[4]),
    .d(al_55bbd6fb),
    .o(al_1dcba582));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~B*~((E*~A))*~(D)+~B*(E*~A)*~(D)+~(~B)*(E*~A)*D+~B*(E*~A)*D))"),
    .INIT(32'h0a0c0f0c))
    al_2375ccfc (
    .a(al_695857c1),
    .b(al_1dcba582),
    .c(al_4002af45),
    .d(al_843f038d),
    .e(al_f65e6902[9]),
    .o(al_8906de47));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fc58ff0d (
    .a(iBusAhb_HRDATA[9]),
    .b(al_b86dd14b[10]),
    .c(al_d518b626),
    .o(al_cf18c1c6[9]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E*~C)*~(F*~(B*~A)))"),
    .INIT(64'h40004400f000ff00))
    al_8d102fa7 (
    .a(al_c7467d2d),
    .b(al_c85e3cfa),
    .c(al_65dc271),
    .d(al_4002af45),
    .e(al_f65e6902[4]),
    .f(al_f65e6902[9]),
    .o(al_9df643fa));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_41b4d49a (
    .a(al_8905c135),
    .b(al_25fbce42[41]),
    .o(al_568af2d5));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(B*~(A*~(~E*~D*~C))))"),
    .INIT(64'hffffffff4444444c))
    al_d445ac77 (
    .a(al_7244a2ec),
    .b(al_52be31ea),
    .c(al_8906de47),
    .d(al_9df643fa),
    .e(al_bdf9a7dd),
    .f(al_568af2d5),
    .o(al_1f3eaa15[9]));
  AL_MAP_LUT6 #(
    .EQN("~(B*~(C)*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+B*C*~((~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))+~(B)*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A)+B*C*(~D*~((~F*~E))*~(A)+~D*(~F*~E)*~(A)+~(~D)*(~F*~E)*A+~D*(~F*~E)*A))"),
    .INIT(64'h3327332733271b0f))
    al_d5478eaa (
    .a(al_bd9d7d67),
    .b(al_cf18c1c6[25]),
    .c(al_cf18c1c6[9]),
    .d(al_a2250ee),
    .e(al_9c16c2f5),
    .f(al_126b3afd[1]),
    .o(al_c524b83f));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_94ad0bd1 (
    .a(al_3629238d),
    .b(al_e2d7fc47),
    .c(al_5fd02584[4]),
    .o(al_f65e6902[4]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_459b532 (
    .a(al_12584de1),
    .b(al_e2d7fc47),
    .c(al_5fd02584[6]),
    .o(al_55bbd6fb));
  AL_MAP_LUT5 #(
    .EQN("~((~B*A)*~((E*~D))*~(C)+(~B*A)*(E*~D)*~(C)+~((~B*A))*(E*~D)*C+(~B*A)*(E*~D)*C)"),
    .INIT(32'hfd0dfdfd))
    al_86f71a62 (
    .a(al_2f34d7b4),
    .b(al_e3502e80),
    .c(al_e2d7fc47),
    .d(al_5fd02584[14]),
    .e(al_5fd02584[15]),
    .o(al_7c8ae043));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~(E*~C)*~(~D*A)))"),
    .INIT(32'h0c8c0088))
    al_746fa90a (
    .a(al_2d6e7982),
    .b(al_3f1d46e5),
    .c(al_a7b01c14[2]),
    .d(al_2c3e73df),
    .e(al_c73c0ba3),
    .o(al_b3684022));
  AL_DFF_X al_8d2f424 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b3684022),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c73c0ba3));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_13a422d5 (
    .a(al_8bea08a7),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[6]),
    .d(al_85a2bdb0[20]),
    .o(al_eb46e9d2));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(~D*C*~B))"),
    .INIT(16'haaba))
    al_3e487ff7 (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[5]),
    .d(al_85a2bdb0[6]),
    .o(al_a8c60ee7));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_8133b89b (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[14]),
    .o(al_9ba628cf));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    al_c234708c (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[13]),
    .d(al_85a2bdb0[14]),
    .o(al_c50e70c2));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_f8d16641 (
    .a(al_8bea08a7),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[6]),
    .o(al_bb2524be));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_f06bd6b4 (
    .a(al_85a2bdb0[3]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[6]),
    .o(al_c52295d9));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~D*~(B*~(~E*~(F*C)))))"),
    .INIT(64'h5544554055445500))
    al_ac0c24be (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[5]),
    .d(al_85a2bdb0[6]),
    .e(al_85a2bdb0[13]),
    .f(al_85a2bdb0[30]),
    .o(al_118827bc));
  AL_MAP_LUT4 #(
    .EQN("(A*~((D*C))*~(B)+A*(D*C)*~(B)+~(A)*(D*C)*B+A*(D*C)*B)"),
    .INIT(16'he222))
    al_450dd54c (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[6]),
    .d(al_85a2bdb0[14]),
    .o(al_4ab1b7b3));
  AL_MAP_LUT4 #(
    .EQN("(A*~((D*B))*~(C)+A*(D*B)*~(C)+~(A)*(D*B)*C+A*(D*B)*C)"),
    .INIT(16'hca0a))
    al_97cb6c0c (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[6]),
    .d(al_85a2bdb0[14]),
    .o(al_40dcfa8c));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    al_af045ffb (
    .a(al_de0f70d9),
    .b(al_85a2bdb0[6]),
    .c(al_85a2bdb0[14]),
    .d(al_85a2bdb0[25]),
    .o(al_361dafb5));
  AL_MAP_LUT6 #(
    .EQN("(E*~D*(A*~((~F*~C))*~(B)+A*(~F*~C)*~(B)+~(A)*(~F*~C)*B+A*(~F*~C)*B))"),
    .INIT(64'h00220000002e0000))
    al_b3895e14 (
    .a(al_85a2bdb0[4]),
    .b(al_85a2bdb0[5]),
    .c(al_85a2bdb0[6]),
    .d(al_85a2bdb0[13]),
    .e(al_85a2bdb0[14]),
    .f(al_85a2bdb0[25]),
    .o(al_c964851));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_16e0c820 (
    .a(al_c964851),
    .b(al_85a2bdb0[2]),
    .c(al_85a2bdb0[12]),
    .o(al_c6966291[20]));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*C*B*~A)"),
    .INIT(64'h0000004000000000))
    al_79346721 (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[5]),
    .d(al_85a2bdb0[6]),
    .e(al_85a2bdb0[14]),
    .f(al_85a2bdb0[25]),
    .o(al_66fb6e33));
  AL_MAP_LUT5 #(
    .EQN("(A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc8c8faf8))
    al_97bc7de8 (
    .a(al_85a2bdb0[5]),
    .b(al_85a2bdb0[6]),
    .c(al_85a2bdb0[14]),
    .d(al_85a2bdb0[25]),
    .e(al_85a2bdb0[30]),
    .o(al_d5b6b580));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*~B*~A)"),
    .INIT(32'h00001000))
    al_5e83a173 (
    .a(al_d5b6b580),
    .b(al_85a2bdb0[2]),
    .c(al_85a2bdb0[4]),
    .d(al_85a2bdb0[12]),
    .e(al_85a2bdb0[13]),
    .o(al_17dd8854));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_4f8914a0 (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[5]),
    .c(al_85a2bdb0[6]),
    .o(al_b8ccdc1c));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_66b4dad (
    .a(al_85a2bdb0[12]),
    .b(al_85a2bdb0[13]),
    .o(al_84a0e6));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*B)*~(C*~A))"),
    .INIT(16'h50dc))
    al_9d333901 (
    .a(al_85a2bdb0[4]),
    .b(al_85a2bdb0[12]),
    .c(al_85a2bdb0[13]),
    .d(al_85a2bdb0[14]),
    .o(al_192b30b5));
  AL_MAP_LUT6 #(
    .EQN("~(~D*~A*(~B*~((F*~E))*~(C)+~B*(F*~E)*~(C)+~(~B)*(F*~E)*C+~B*(F*~E)*C))"),
    .INIT(64'hfffeffaefffefffe))
    al_9a56fa9e (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[5]),
    .d(al_85a2bdb0[6]),
    .e(al_85a2bdb0[14]),
    .f(al_85a2bdb0[25]),
    .o(al_4a753b95[11]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h222200222e2e00ee))
    al_9c13ee16 (
    .a(al_85a2bdb0[4]),
    .b(al_85a2bdb0[5]),
    .c(al_85a2bdb0[6]),
    .d(al_85a2bdb0[12]),
    .e(al_85a2bdb0[13]),
    .f(al_85a2bdb0[25]),
    .o(al_acac884e));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_65f67d3c (
    .a(al_acac884e),
    .b(al_85a2bdb0[2]),
    .o(al_c0c7b1b4));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    al_62e1487a (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_98804c07),
    .d(al_bf952132),
    .o(al_6e268dd3[10]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    al_6293a57d (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_3ebb68c3),
    .d(al_76a52f3d),
    .o(al_6e268dd3[11]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    al_829e9f32 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_d00a6f56),
    .d(al_c861c8f0),
    .o(al_6e268dd3[12]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    al_29bdbb86 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_e6455839),
    .d(al_8a841cb4),
    .o(al_6e268dd3[13]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    al_9a91c891 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_7e6320f4),
    .d(al_33a2911e),
    .o(al_6e268dd3[14]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    al_7686cbce (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_f61ec828),
    .d(al_73fb1ee5),
    .o(al_6e268dd3[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3dcde852 (
    .a(dBusAhb_HSIZE[1]),
    .b(al_7d27d680),
    .c(al_f4b5275b),
    .o(al_6e268dd3[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_395ebb09 (
    .a(dBusAhb_HSIZE[1]),
    .b(al_d76255c5),
    .c(al_2370214),
    .o(al_6e268dd3[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d72f5bf (
    .a(dBusAhb_HSIZE[1]),
    .b(al_3b0f4da7),
    .c(al_bf952132),
    .o(al_6e268dd3[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bb9cc356 (
    .a(dBusAhb_HSIZE[1]),
    .b(al_c7df4b4d),
    .c(al_76a52f3d),
    .o(al_6e268dd3[19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d989661b (
    .a(dBusAhb_HSIZE[1]),
    .b(al_a831c176),
    .c(al_c861c8f0),
    .o(al_6e268dd3[20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f184a9bb (
    .a(dBusAhb_HSIZE[1]),
    .b(al_658bb789),
    .c(al_8a841cb4),
    .o(al_6e268dd3[21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_34b9ac7f (
    .a(dBusAhb_HSIZE[1]),
    .b(al_ffc4fe26),
    .c(al_33a2911e),
    .o(al_6e268dd3[22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_585a0977 (
    .a(dBusAhb_HSIZE[1]),
    .b(al_1f5093b5),
    .c(al_73fb1ee5),
    .o(al_6e268dd3[23]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_a2e1f044 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_53b3dbc6),
    .d(al_bdb28b76),
    .e(al_f4b5275b),
    .o(al_6e268dd3[24]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_dbae8965 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_e611ec68),
    .d(al_6d92b3c6),
    .e(al_2370214),
    .o(al_6e268dd3[25]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_831009c6 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_6ec45564),
    .d(al_98804c07),
    .e(al_bf952132),
    .o(al_6e268dd3[26]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_2c47cf93 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_102b7ad2),
    .d(al_3ebb68c3),
    .e(al_76a52f3d),
    .o(al_6e268dd3[27]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_cb0ea20e (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_3b8c31d7),
    .d(al_d00a6f56),
    .e(al_c861c8f0),
    .o(al_6e268dd3[28]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_4d9dca7 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_3626cb0),
    .d(al_e6455839),
    .e(al_8a841cb4),
    .o(al_6e268dd3[29]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_8bc53604 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_f1bb92e9),
    .d(al_7e6320f4),
    .e(al_33a2911e),
    .o(al_6e268dd3[30]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_a9f4a66b (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_60dd36d7),
    .d(al_f61ec828),
    .e(al_73fb1ee5),
    .o(al_6e268dd3[31]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    al_36212611 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_bdb28b76),
    .d(al_f4b5275b),
    .o(al_6e268dd3[8]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    al_3fabd927 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_6d92b3c6),
    .d(al_2370214),
    .o(al_6e268dd3[9]));
  AL_MAP_LUT5 #(
    .EQN("(C*~((~E*~D*A))*~(B)+C*(~E*~D*A)*~(B)+~(C)*(~E*~D*A)*B+C*(~E*~D*A)*B)"),
    .INIT(32'h303030b8))
    al_ea6aceed (
    .a(al_1a09507b),
    .b(dBusAhb_HREADY_IN),
    .c(al_d020f13b),
    .d(al_b8fe1a1f),
    .e(dBusAhb_HWRITE),
    .o(al_3d9557e1));
  AL_DFF_X al_b6afdbff (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3d9557e1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d020f13b));
  AL_MAP_LUT6 #(
    .EQN("(C*B*A*~(D*~(E)*~(F)+D*E*~(F)+~(D)*E*F+D*E*F))"),
    .INIT(64'h0000808000800080))
    al_85340105 (
    .a(al_8bea08a7),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[6]),
    .d(al_85a2bdb0[20]),
    .e(al_85a2bdb0[21]),
    .f(al_85a2bdb0[28]),
    .o(al_40a6f08c[27]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf5a0f5a0dddd8888))
    al_1ea49ce3 (
    .a(al_f2330f79[0]),
    .b(al_18077581[2]),
    .c(al_18077581[29]),
    .d(al_18077581[28]),
    .e(al_18077581[3]),
    .f(al_a994b7f),
    .o(al_660ff49e));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_dd1fc344 (
    .a(al_5d89de3c),
    .b(al_7428b0ee),
    .c(al_f2330f79[2]),
    .o(al_1fb1fe24));
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(D)*~(E)+C*D*~(E)+~(C)*D*E+C*D*E))*~(B)+A*(C*~(D)*~(E)+C*D*~(E)+~(C)*D*E+C*D*E)*~(B)+~(A)*(C*~(D)*~(E)+C*D*~(E)+~(C)*D*E+C*D*E)*B+A*(C*~(D)*~(E)+C*D*~(E)+~(C)*D*E+C*D*E)*B)"),
    .INIT(32'hee22e2e2))
    al_a0cc062e (
    .a(al_660ff49e),
    .b(al_f2330f79[1]),
    .c(al_18077581[1]),
    .d(al_18077581[30]),
    .e(al_a994b7f),
    .o(al_5a1a38b6));
  AL_MAP_LUT6 #(
    .EQN("~(A*~((E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F))*~((C*B))+A*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*~((C*B))+~(A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*(C*B)+A*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*(C*B))"),
    .INIT(64'h15d515d51515d5d5))
    al_6b7b0626 (
    .a(al_5a1a38b6),
    .b(al_f2330f79[1]),
    .c(al_f2330f79[0]),
    .d(al_18077581[31]),
    .e(al_18077581[0]),
    .f(al_a994b7f),
    .o(al_2b49ac1e));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f00ff3333aaaa))
    al_af34c066 (
    .a(al_13f338be),
    .b(al_1fb1fe24),
    .c(al_2b49ac1e),
    .d(al_e9d7a836),
    .e(al_786d2b97),
    .f(al_ea114973),
    .o(al_9e82589f[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h3333f0f05555ff00))
    al_2d024325 (
    .a(al_71df23fe),
    .b(al_8953e749),
    .c(al_87fbe8d),
    .d(al_ee1342f7[32]),
    .e(al_f2330f79[4]),
    .f(al_f2330f79[3]),
    .o(al_9e82589f[10]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_d31a3a61 (
    .a(al_48e8a022),
    .b(al_c21c784f),
    .c(al_f2330f79[2]),
    .o(al_de36fb50));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_7a9baf70 (
    .a(al_271d0926),
    .b(al_ac27d20b),
    .c(al_f2330f79[2]),
    .o(al_4f8cbab6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h333355550f0fff00))
    al_25c610ba (
    .a(al_4381d4c9),
    .b(al_4f8cbab6),
    .c(al_de36fb50),
    .d(al_ee1342f7[32]),
    .e(al_f2330f79[4]),
    .f(al_f2330f79[3]),
    .o(al_9e82589f[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h3333aaaa0f0fff00))
    al_f0e24c93 (
    .a(al_bdd9239c),
    .b(al_d1b00369),
    .c(al_a4f54b87),
    .d(al_ee1342f7[32]),
    .e(al_f2330f79[4]),
    .f(al_f2330f79[3]),
    .o(al_9e82589f[12]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_86763e72 (
    .a(al_ac17e182),
    .b(al_74831af1),
    .c(al_f2330f79[1]),
    .o(al_99df9c8d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h3333aaaa0f0fff00))
    al_7f295810 (
    .a(al_d14a1180),
    .b(al_efb93bad),
    .c(al_897eb9f3),
    .d(al_ee1342f7[32]),
    .e(al_f2330f79[4]),
    .f(al_f2330f79[3]),
    .o(al_9e82589f[13]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_5307e1fa (
    .a(al_97966a28),
    .b(al_ae1d4fee),
    .c(al_f2330f79[1]),
    .o(al_470c29ce));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_aa80172e (
    .a(al_5281bd0f),
    .b(al_784638ef),
    .c(al_f2330f79[1]),
    .o(al_7ba3de08));
  AL_MAP_LUT6 #(
    .EQN("(~(D*~(E)*~((F@C))+D*E*~((F@C))+~(D)*E*(F@C)+D*E*(F@C))*~(A)*~(B)+~(D*~(E)*~((F@C))+D*E*~((F@C))+~(D)*E*(F@C)+D*E*(F@C))*A*~(B)+~(~(D*~(E)*~((F@C))+D*E*~((F@C))+~(D)*E*(F@C)+D*E*(F@C)))*A*B+~(D*~(E)*~((F@C))+D*E*~((F@C))+~(D)*E*(F@C)+D*E*(F@C))*A*B)"),
    .INIT(64'h88b88bbb888bb8bb))
    al_5a7711ab (
    .a(al_723a595b),
    .b(al_f2330f79[1]),
    .c(al_f2330f79[0]),
    .d(al_18077581[16]),
    .e(al_18077581[15]),
    .f(al_a994b7f),
    .o(al_6c7e2f3));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_4104aedc (
    .a(al_99df9c8d),
    .b(al_7ba3de08),
    .c(al_f2330f79[2]),
    .o(al_897eb9f3));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    al_7565506f (
    .a(al_6c7e2f3),
    .b(al_470c29ce),
    .c(al_f2330f79[2]),
    .o(al_efb93bad));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D*C))+A*B*~((D*C))+~(A)*B*(D*C)+A*B*(D*C))"),
    .INIT(16'h3555))
    al_d30257 (
    .a(al_ee1342f7[32]),
    .b(al_6d9a66ce),
    .c(al_3789ddb5),
    .d(al_f2330f79[1]),
    .o(al_fc3546f));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_e248e68 (
    .a(al_a7eb7455),
    .b(al_9ba605ab),
    .c(al_f2330f79[2]),
    .o(al_c14f8945));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_3676503d (
    .a(al_1b1495c6),
    .b(al_39f4f94a),
    .c(al_f2330f79[2]),
    .o(al_3a175d67));
  AL_MAP_LUT5 #(
    .EQN("~(C*~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*~(D)+C*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(D)+~(C)*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*D+C*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*D)"),
    .INIT(32'h330f550f))
    al_79cdc51b (
    .a(al_c14f8945),
    .b(al_3a175d67),
    .c(al_fc3546f),
    .d(al_f2330f79[4]),
    .e(al_f2330f79[3]),
    .o(al_9e82589f[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'he4e4e4e4ffaa5500))
    al_30bdba85 (
    .a(al_f2330f79[0]),
    .b(al_18077581[1]),
    .c(al_18077581[2]),
    .d(al_18077581[30]),
    .e(al_18077581[29]),
    .f(al_a994b7f),
    .o(al_28aac2f6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F)"),
    .INIT(64'h0055aaff1b1b1b1b))
    al_3a5c6fb6 (
    .a(al_f2330f79[0]),
    .b(al_18077581[22]),
    .c(al_18077581[21]),
    .d(al_18077581[9]),
    .e(al_18077581[10]),
    .f(al_a994b7f),
    .o(al_784638ef));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_1e456618 (
    .a(al_28aac2f6),
    .b(al_ac17e182),
    .c(al_f2330f79[1]),
    .o(al_8bfeeae9));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_35984ec2 (
    .a(al_ae1d4fee),
    .b(al_784638ef),
    .c(al_f2330f79[1]),
    .o(al_48e8a022));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_c28dffaf (
    .a(al_74831af1),
    .b(al_5281bd0f),
    .c(al_f2330f79[1]),
    .o(al_c21c784f));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((D*~(E)*~((F@C))+D*E*~((F@C))+~(D)*E*(F@C)+D*E*(F@C)))*~(B)+~A*(D*~(E)*~((F@C))+D*E*~((F@C))+~(D)*E*(F@C)+D*E*(F@C))*~(B)+~(~A)*(D*~(E)*~((F@C))+D*E*~((F@C))+~(D)*E*(F@C)+D*E*(F@C))*B+~A*(D*~(E)*~((F@C))+D*E*~((F@C))+~(D)*E*(F@C)+D*E*(F@C))*B)"),
    .INIT(64'hdd1dd111ddd11d11))
    al_e654742b (
    .a(al_97966a28),
    .b(al_f2330f79[1]),
    .c(al_f2330f79[0]),
    .d(al_18077581[16]),
    .e(al_18077581[15]),
    .f(al_a994b7f),
    .o(al_271d0926));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_432e79ce (
    .a(al_8bfeeae9),
    .b(al_c21c784f),
    .c(al_f2330f79[2]),
    .o(al_f6c0774b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff55aa00e4e4e4e4))
    al_91a13de6 (
    .a(al_f2330f79[0]),
    .b(al_18077581[28]),
    .c(al_18077581[27]),
    .d(al_18077581[4]),
    .e(al_18077581[3]),
    .f(al_a994b7f),
    .o(al_ac17e182));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_f859630b (
    .a(al_271d0926),
    .b(al_48e8a022),
    .c(al_f2330f79[2]),
    .o(al_3833a138));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h5555fff03333f0f0))
    al_ea8a3fff (
    .a(al_3833a138),
    .b(al_f6c0774b),
    .c(al_ee1342f7[32]),
    .d(al_2dba6136),
    .e(al_f2330f79[4]),
    .f(al_f2330f79[3]),
    .o(al_9e82589f[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F)"),
    .INIT(64'h0055aaff1b1b1b1b))
    al_80a62c40 (
    .a(al_f2330f79[0]),
    .b(al_18077581[26]),
    .c(al_18077581[25]),
    .d(al_18077581[5]),
    .e(al_18077581[6]),
    .f(al_a994b7f),
    .o(al_74831af1));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00aa55ff1b1b1b1b))
    al_99c931ce (
    .a(al_f2330f79[0]),
    .b(al_18077581[18]),
    .c(al_18077581[17]),
    .d(al_18077581[14]),
    .e(al_18077581[13]),
    .f(al_a994b7f),
    .o(al_97966a28));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00aa55ff1b1b1b1b))
    al_435dd5d4 (
    .a(al_f2330f79[0]),
    .b(al_18077581[20]),
    .c(al_18077581[19]),
    .d(al_18077581[12]),
    .e(al_18077581[11]),
    .f(al_a994b7f),
    .o(al_ae1d4fee));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F)"),
    .INIT(64'h0055aaff1b1b1b1b))
    al_511bf588 (
    .a(al_f2330f79[0]),
    .b(al_18077581[24]),
    .c(al_18077581[23]),
    .d(al_18077581[7]),
    .e(al_18077581[8]),
    .f(al_a994b7f),
    .o(al_5281bd0f));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_8a7d1cd0 (
    .a(al_d9533dba),
    .b(al_5b8651b5),
    .c(al_f2330f79[2]),
    .o(al_d9a23597));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_5b52cb2 (
    .a(al_f9c1044d),
    .b(al_69c28a29),
    .c(al_f2330f79[2]),
    .o(al_76cdacda));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_90d817fa (
    .a(al_d9a23597),
    .b(al_76cdacda),
    .c(al_f2330f79[3]),
    .o(al_13f338be));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_597e060d (
    .a(al_13f338be),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[16]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_ac0f756b (
    .a(al_3c39e4b0),
    .b(al_3c3c44e5),
    .c(al_f2330f79[3]),
    .o(al_7b0b987));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_aafcc084 (
    .a(al_7b0b987),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[17]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_35373447 (
    .a(al_951b8fda),
    .b(al_a7a12e87),
    .c(al_f2330f79[1]),
    .o(al_a7eb7455));
  AL_MAP_LUT5 #(
    .EQN("((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haaf0aacc))
    al_812ac476 (
    .a(al_a7eb7455),
    .b(al_ee1342f7[32]),
    .c(al_6d9a66ce),
    .d(al_f2330f79[2]),
    .e(al_f2330f79[1]),
    .o(al_87fbe8d));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_1ccf6c07 (
    .a(al_7daf0c48),
    .b(al_fb6b4008),
    .c(al_f2330f79[1]),
    .o(al_9ba605ab));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_54a7899f (
    .a(al_18e8ea79),
    .b(al_d41aa0e7),
    .c(al_f2330f79[1]),
    .o(al_39f4f94a));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_45218a0b (
    .a(al_9ba605ab),
    .b(al_39f4f94a),
    .c(al_f2330f79[2]),
    .o(al_71df23fe));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_11f07d59 (
    .a(al_71df23fe),
    .b(al_87fbe8d),
    .c(al_f2330f79[3]),
    .o(al_fb1aae));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a5835075 (
    .a(al_fb1aae),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[18]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_91510d4b (
    .a(al_4381d4c9),
    .b(al_de36fb50),
    .c(al_f2330f79[3]),
    .o(al_b8cddd4));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_46f1f1f1 (
    .a(al_b8cddd4),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[19]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf0f0aaaaff00cccc))
    al_adeb1ece (
    .a(al_18077581[1]),
    .b(al_18077581[2]),
    .c(al_18077581[30]),
    .d(al_18077581[29]),
    .e(al_a994b7f),
    .f(al_f2330f79[0]),
    .o(al_68a3d338));
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'hccaaf0aa))
    al_6a64a270 (
    .a(al_20e2d49e),
    .b(al_68a3d338),
    .c(al_2c5a98b1),
    .d(al_f2330f79[2]),
    .e(al_f2330f79[1]),
    .o(al_8a026941));
  AL_MAP_LUT5 #(
    .EQN("(A*~((~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E))*~(D)+A*(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*~(D)+~(A)*(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*D+A*(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*D)"),
    .INIT(32'hf0aa33aa))
    al_fc35bad9 (
    .a(al_7b0b987),
    .b(al_2edab7d3),
    .c(al_8a026941),
    .d(al_f2330f79[4]),
    .e(al_f2330f79[3]),
    .o(al_9e82589f[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E))*~(B)+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*~(B)+~(~A)*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)"),
    .INIT(32'hd1d1dd11))
    al_46c2c0f (
    .a(al_4e9ff654),
    .b(al_f2330f79[0]),
    .c(al_18077581[1]),
    .d(al_18077581[30]),
    .e(al_a994b7f),
    .o(al_6d9a66ce));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_d9ed4feb (
    .a(al_a7a12e87),
    .b(al_7daf0c48),
    .c(al_f2330f79[1]),
    .o(al_5b8651b5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F)"),
    .INIT(64'h0055aaff1b1b1b1b))
    al_c20d4590 (
    .a(al_f2330f79[0]),
    .b(al_18077581[23]),
    .c(al_18077581[22]),
    .d(al_18077581[8]),
    .e(al_18077581[9]),
    .f(al_a994b7f),
    .o(al_fb6b4008));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F)"),
    .INIT(64'h0055aaff1b1b1b1b))
    al_4503b9ab (
    .a(al_f2330f79[0]),
    .b(al_18077581[21]),
    .c(al_18077581[20]),
    .d(al_18077581[10]),
    .e(al_18077581[11]),
    .f(al_a994b7f),
    .o(al_d41aa0e7));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_9bd233eb (
    .a(al_fb6b4008),
    .b(al_d41aa0e7),
    .c(al_f2330f79[1]),
    .o(al_69c28a29));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_165aec3d (
    .a(al_5b8651b5),
    .b(al_69c28a29),
    .c(al_f2330f79[2]),
    .o(al_a4f54b87));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_f1e0fbc6 (
    .a(al_bdd9239c),
    .b(al_a4f54b87),
    .c(al_f2330f79[3]),
    .o(al_2d4bf1ba));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8be908a7 (
    .a(al_2d4bf1ba),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[20]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeee4444fa50fa50))
    al_18c68842 (
    .a(al_f2330f79[0]),
    .b(al_18077581[2]),
    .c(al_18077581[29]),
    .d(al_18077581[28]),
    .e(al_18077581[3]),
    .f(al_a994b7f),
    .o(al_951b8fda));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_cb9c075c (
    .a(al_6d9a66ce),
    .b(al_951b8fda),
    .c(al_f2330f79[1]),
    .o(al_d9533dba));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_5725bbfd (
    .a(al_d9533dba),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[2]),
    .o(al_bdd9239c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F)"),
    .INIT(64'h0055aaff1b1b1b1b))
    al_e1e599e7 (
    .a(al_f2330f79[0]),
    .b(al_18077581[27]),
    .c(al_18077581[26]),
    .d(al_18077581[4]),
    .e(al_18077581[5]),
    .f(al_a994b7f),
    .o(al_a7a12e87));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F)"),
    .INIT(64'h0055aaff1b1b1b1b))
    al_58e1ce3d (
    .a(al_f2330f79[0]),
    .b(al_18077581[25]),
    .c(al_18077581[24]),
    .d(al_18077581[6]),
    .e(al_18077581[7]),
    .f(al_a994b7f),
    .o(al_7daf0c48));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_fcfacafa (
    .a(al_d14a1180),
    .b(al_897eb9f3),
    .c(al_f2330f79[3]),
    .o(al_a840afb1));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_dd6a9882 (
    .a(al_a840afb1),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_37c0721f (
    .a(al_220ba3d7),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[22]));
  AL_MAP_LUT4 #(
    .EQN("~((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D)"),
    .INIT(16'h55fc))
    al_743ace5b (
    .a(al_f6c0774b),
    .b(al_ee1342f7[32]),
    .c(al_2dba6136),
    .d(al_f2330f79[3]),
    .o(al_95cc331e));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_456a7e62 (
    .a(al_95cc331e),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[23]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_c5b2127d (
    .a(al_d9a23597),
    .b(al_ee1342f7[32]),
    .c(al_ea114973),
    .o(al_9e82589f[24]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_13cb58ed (
    .a(al_4cc73535),
    .b(al_99df9c8d),
    .c(al_f2330f79[2]),
    .o(al_3c39e4b0));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_e7f8fff9 (
    .a(al_3c39e4b0),
    .b(al_ee1342f7[32]),
    .c(al_ea114973),
    .o(al_9e82589f[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2049d0e1 (
    .a(al_87fbe8d),
    .b(al_ee1342f7[32]),
    .c(al_ea114973),
    .o(al_9e82589f[26]));
  AL_MAP_LUT6 #(
    .EQN("((~B*~(F*E*~C))*~(A)*~(D)+(~B*~(F*E*~C))*A*~(D)+~((~B*~(F*E*~C)))*A*D+(~B*~(F*E*~C))*A*D)"),
    .INIT(64'haa30aa33aa33aa33))
    al_10263a3f (
    .a(al_8bfeeae9),
    .b(al_ee1342f7[32]),
    .c(al_4e9ff654),
    .d(al_f2330f79[2]),
    .e(al_f2330f79[1]),
    .f(al_f2330f79[0]),
    .o(al_4381d4c9));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_6fd34ea4 (
    .a(al_4381d4c9),
    .b(al_ee1342f7[32]),
    .c(al_ea114973),
    .o(al_9e82589f[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2b15a95c (
    .a(al_bdd9239c),
    .b(al_ee1342f7[32]),
    .c(al_ea114973),
    .o(al_9e82589f[28]));
  AL_MAP_LUT5 #(
    .EQN("~(~(~A*~(E*~C))*~(B)*~(D)+~(~A*~(E*~C))*B*~(D)+~(~(~A*~(E*~C)))*B*D+~(~A*~(E*~C))*B*D)"),
    .INIT(32'h33503355))
    al_adb97ef2 (
    .a(al_ee1342f7[32]),
    .b(al_28aac2f6),
    .c(al_4e9ff654),
    .d(al_f2330f79[1]),
    .e(al_f2330f79[0]),
    .o(al_4cc73535));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_2e595de0 (
    .a(al_4cc73535),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[2]),
    .o(al_d14a1180));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_faddd172 (
    .a(al_d14a1180),
    .b(al_ee1342f7[32]),
    .c(al_ea114973),
    .o(al_9e82589f[29]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_5371bdf9 (
    .a(al_be8dbeba),
    .b(al_460aa351),
    .c(al_f2330f79[1]),
    .o(al_1b1495c6));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_45f3c5df (
    .a(al_4183cccb),
    .b(al_f405df5e),
    .c(al_f2330f79[1]),
    .o(al_e92fad27));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_c7b69186 (
    .a(al_cb204385),
    .b(al_fb048e7c),
    .c(al_f2330f79[1]),
    .o(al_8f3d3123));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_47b8a68d (
    .a(al_1b1495c6),
    .b(al_8f3d3123),
    .c(al_f2330f79[2]),
    .o(al_8953e749));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0033aa0fff33aa))
    al_10832ccc (
    .a(al_8953e749),
    .b(al_e92fad27),
    .c(al_660ff49e),
    .d(al_30a65d08),
    .e(al_3789ddb5),
    .f(al_5824822d),
    .o(al_6c0635b4));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_69d2d891 (
    .a(al_fb1aae),
    .b(al_6c0635b4),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[2]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_c1d3bc97 (
    .a(al_fc3546f),
    .b(al_ee1342f7[32]),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[30]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_849ea145 (
    .a(al_27c2eb8[0]),
    .b(al_27c2eb8[1]),
    .o(al_a994b7f));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_6bd8d3c2 (
    .a(al_18077581[31]),
    .b(al_18077581[0]),
    .c(al_a994b7f),
    .o(al_4e9ff654));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_c525e52a (
    .a(al_4e9ff654),
    .b(al_27c2eb8[0]),
    .c(al_27c2eb8[1]),
    .o(al_ee1342f7[32]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_1ac2ce5f (
    .a(al_f2330f79[4]),
    .b(al_f2330f79[3]),
    .o(al_ea114973));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    al_24de9c77 (
    .a(al_4e9ff654),
    .b(al_f2330f79[2]),
    .c(al_f2330f79[1]),
    .d(al_f2330f79[0]),
    .o(al_2dba6136));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    al_1ebe6c46 (
    .a(al_ee1342f7[32]),
    .b(al_2dba6136),
    .c(al_ea114973),
    .o(al_9e82589f[31]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_5fdfc3f (
    .a(al_f2330f79[3]),
    .b(al_f2330f79[2]),
    .o(al_3789ddb5));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_790a06ac (
    .a(al_b8cddd4),
    .b(al_cf16e2e3),
    .c(al_f2330f79[4]),
    .o(al_9e82589f[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    al_1c7b1994 (
    .a(al_f2330f79[3]),
    .b(al_f2330f79[2]),
    .c(al_f2330f79[1]),
    .o(al_30a65d08));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h2727272700aa55ff))
    al_7353a3f3 (
    .a(al_f2330f79[0]),
    .b(al_18077581[26]),
    .c(al_18077581[25]),
    .d(al_18077581[5]),
    .e(al_18077581[6]),
    .f(al_a994b7f),
    .o(al_9617ef5a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hd8d8d8d8ffaa5500))
    al_2b7a7a7c (
    .a(al_f2330f79[0]),
    .b(al_18077581[28]),
    .c(al_18077581[27]),
    .d(al_18077581[4]),
    .e(al_18077581[3]),
    .f(al_a994b7f),
    .o(al_2c5a98b1));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0fff33aa0f0033aa))
    al_3835de17 (
    .a(al_4f8cbab6),
    .b(al_61365560),
    .c(al_2c5a98b1),
    .d(al_30a65d08),
    .e(al_3789ddb5),
    .f(al_9617ef5a),
    .o(al_cf16e2e3));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00aa55ff1b1b1b1b))
    al_e2c21d60 (
    .a(al_f2330f79[0]),
    .b(al_18077581[17]),
    .c(al_18077581[16]),
    .d(al_18077581[15]),
    .e(al_18077581[14]),
    .f(al_a994b7f),
    .o(al_be8dbeba));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h272727270055aaff))
    al_a00d61d6 (
    .a(al_f2330f79[0]),
    .b(al_18077581[19]),
    .c(al_18077581[18]),
    .d(al_18077581[13]),
    .e(al_18077581[12]),
    .f(al_a994b7f),
    .o(al_cb204385));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h2727272700aa55ff))
    al_a21a0608 (
    .a(al_f2330f79[0]),
    .b(al_18077581[21]),
    .c(al_18077581[20]),
    .d(al_18077581[10]),
    .e(al_18077581[11]),
    .f(al_a994b7f),
    .o(al_fb048e7c));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hd8d8d8d8ff55aa00))
    al_29dc3756 (
    .a(al_f2330f79[0]),
    .b(al_18077581[27]),
    .c(al_18077581[26]),
    .d(al_18077581[4]),
    .e(al_18077581[5]),
    .f(al_a994b7f),
    .o(al_5824822d));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_6ac01567 (
    .a(al_18e8ea79),
    .b(al_be8dbeba),
    .c(al_f2330f79[1]),
    .o(al_f9c1044d));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_2dd058fe (
    .a(al_460aa351),
    .b(al_cb204385),
    .c(al_f2330f79[1]),
    .o(al_5d89de3c));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_5763cd50 (
    .a(al_4183cccb),
    .b(al_fb048e7c),
    .c(al_f2330f79[1]),
    .o(al_7428b0ee));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_5db31d69 (
    .a(al_f405df5e),
    .b(al_5824822d),
    .c(al_f2330f79[1]),
    .o(al_e9d7a836));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_d93378d7 (
    .a(al_f9c1044d),
    .b(al_5d89de3c),
    .c(al_f2330f79[2]),
    .o(al_d1b00369));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00fff0f03333aaaa))
    al_ecfd76db (
    .a(al_2d4bf1ba),
    .b(al_d1b00369),
    .c(al_7428b0ee),
    .d(al_e9d7a836),
    .e(al_786d2b97),
    .f(al_ea114973),
    .o(al_9e82589f[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h272727270055aaff))
    al_d8ff8036 (
    .a(al_f2330f79[0]),
    .b(al_18077581[17]),
    .c(al_18077581[16]),
    .d(al_18077581[15]),
    .e(al_18077581[14]),
    .f(al_a994b7f),
    .o(al_460aa351));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00aa55ff1b1b1b1b))
    al_557121e2 (
    .a(al_f2330f79[0]),
    .b(al_18077581[19]),
    .c(al_18077581[18]),
    .d(al_18077581[13]),
    .e(al_18077581[12]),
    .f(al_a994b7f),
    .o(al_18e8ea79));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h2727272700aa55ff))
    al_15a24c67 (
    .a(al_f2330f79[0]),
    .b(al_18077581[23]),
    .c(al_18077581[22]),
    .d(al_18077581[8]),
    .e(al_18077581[9]),
    .f(al_a994b7f),
    .o(al_4183cccb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h2727272700aa55ff))
    al_6fe43e40 (
    .a(al_f2330f79[0]),
    .b(al_18077581[25]),
    .c(al_18077581[24]),
    .d(al_18077581[6]),
    .e(al_18077581[7]),
    .f(al_a994b7f),
    .o(al_f405df5e));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_24fceb67 (
    .a(al_42c07e1a),
    .b(al_d6c2acee),
    .c(al_f2330f79[1]),
    .o(al_5fe9efd2));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_dee5582c (
    .a(al_dd28d822),
    .b(al_9617ef5a),
    .c(al_f2330f79[1]),
    .o(al_20e2d49e));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf0f0ff003333aaaa))
    al_25cdc1ba (
    .a(al_a840afb1),
    .b(al_efb93bad),
    .c(al_20e2d49e),
    .d(al_5fe9efd2),
    .e(al_786d2b97),
    .f(al_ea114973),
    .o(al_9e82589f[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(B*~(C)*~((F*E))+B*C*~((F*E))+~(B)*C*(F*E)+B*C*(F*E))*~(A)*~(D)+~(B*~(C)*~((F*E))+B*C*~((F*E))+~(B)*C*(F*E)+B*C*(F*E))*A*~(D)+~(~(B*~(C)*~((F*E))+B*C*~((F*E))+~(B)*C*(F*E)+B*C*(F*E)))*A*D+~(B*~(C)*~((F*E))+B*C*~((F*E))+~(B)*C*(F*E)+B*C*(F*E))*A*D)"),
    .INIT(64'h55f055cc55cc55cc))
    al_bee1d804 (
    .a(al_c14f8945),
    .b(al_ee1342f7[32]),
    .c(al_6d9a66ce),
    .d(al_f2330f79[3]),
    .e(al_f2330f79[2]),
    .f(al_f2330f79[1]),
    .o(al_220ba3d7));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf0f0ff003333aaaa))
    al_c7cacd75 (
    .a(al_220ba3d7),
    .b(al_3a175d67),
    .c(al_e92fad27),
    .d(al_8f3d3123),
    .e(al_786d2b97),
    .f(al_ea114973),
    .o(al_9e82589f[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    al_646c7677 (
    .a(al_f2330f79[4]),
    .b(al_f2330f79[3]),
    .c(al_f2330f79[2]),
    .o(al_786d2b97));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_3308699 (
    .a(al_723a595b),
    .b(al_42c07e1a),
    .c(al_f2330f79[1]),
    .o(al_ac27d20b));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_f577a18c (
    .a(al_dd28d822),
    .b(al_d6c2acee),
    .c(al_f2330f79[1]),
    .o(al_61365560));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf0f0ff003333aaaa))
    al_b907b3e5 (
    .a(al_95cc331e),
    .b(al_3833a138),
    .c(al_61365560),
    .d(al_ac27d20b),
    .e(al_786d2b97),
    .f(al_ea114973),
    .o(al_9e82589f[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h272727270055aaff))
    al_df62cad6 (
    .a(al_f2330f79[0]),
    .b(al_18077581[18]),
    .c(al_18077581[17]),
    .d(al_18077581[14]),
    .e(al_18077581[13]),
    .f(al_a994b7f),
    .o(al_723a595b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h272727270055aaff))
    al_89e2cdba (
    .a(al_f2330f79[0]),
    .b(al_18077581[20]),
    .c(al_18077581[19]),
    .d(al_18077581[12]),
    .e(al_18077581[11]),
    .f(al_a994b7f),
    .o(al_42c07e1a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h2727272700aa55ff))
    al_e96a191d (
    .a(al_f2330f79[0]),
    .b(al_18077581[22]),
    .c(al_18077581[21]),
    .d(al_18077581[9]),
    .e(al_18077581[10]),
    .f(al_a994b7f),
    .o(al_d6c2acee));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h2727272700aa55ff))
    al_f81013ef (
    .a(al_f2330f79[0]),
    .b(al_18077581[24]),
    .c(al_18077581[23]),
    .d(al_18077581[7]),
    .e(al_18077581[8]),
    .f(al_a994b7f),
    .o(al_dd28d822));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f0f55553333ff00))
    al_1863f9bd (
    .a(al_d9a23597),
    .b(al_76cdacda),
    .c(al_1fb1fe24),
    .d(al_ee1342f7[32]),
    .e(al_f2330f79[4]),
    .f(al_f2330f79[3]),
    .o(al_9e82589f[8]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_21d05144 (
    .a(al_470c29ce),
    .b(al_7ba3de08),
    .c(al_f2330f79[2]),
    .o(al_3c3c44e5));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_eaf29ce7 (
    .a(al_6c7e2f3),
    .b(al_5fe9efd2),
    .c(al_f2330f79[2]),
    .o(al_2edab7d3));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h333355550f0fff00))
    al_274a812a (
    .a(al_3c39e4b0),
    .b(al_2edab7d3),
    .c(al_3c3c44e5),
    .d(al_ee1342f7[32]),
    .e(al_f2330f79[4]),
    .f(al_f2330f79[3]),
    .o(al_9e82589f[9]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_5a61b914 (
    .a(al_f2330f79[0]),
    .b(al_df7b4407),
    .o(al_3ca44efd[0]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_2bc0e599 (
    .a(al_f2330f79[10]),
    .b(al_df7b4407),
    .o(al_3ca44efd[10]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_2b8f0569 (
    .a(al_f2330f79[11]),
    .b(al_df7b4407),
    .o(al_3ca44efd[11]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_b43fd421 (
    .a(al_f2330f79[12]),
    .b(al_df7b4407),
    .o(al_3ca44efd[12]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_6d0f7d8b (
    .a(al_f2330f79[13]),
    .b(al_df7b4407),
    .o(al_3ca44efd[13]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_27d93c4a (
    .a(al_f2330f79[14]),
    .b(al_df7b4407),
    .o(al_3ca44efd[14]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_51998e5c (
    .a(al_f2330f79[15]),
    .b(al_df7b4407),
    .o(al_3ca44efd[15]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_1937f971 (
    .a(al_f2330f79[16]),
    .b(al_df7b4407),
    .o(al_3ca44efd[16]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_a474b9b2 (
    .a(al_f2330f79[17]),
    .b(al_df7b4407),
    .o(al_3ca44efd[17]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_9929930 (
    .a(al_f2330f79[18]),
    .b(al_df7b4407),
    .o(al_3ca44efd[18]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_bf872c9a (
    .a(al_f2330f79[19]),
    .b(al_df7b4407),
    .o(al_3ca44efd[19]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_8c2f7daf (
    .a(al_f2330f79[1]),
    .b(al_df7b4407),
    .o(al_3ca44efd[1]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_be328864 (
    .a(al_f2330f79[20]),
    .b(al_df7b4407),
    .o(al_3ca44efd[20]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_4a228c5c (
    .a(al_f2330f79[21]),
    .b(al_df7b4407),
    .o(al_3ca44efd[21]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_9c8931ed (
    .a(al_f2330f79[22]),
    .b(al_df7b4407),
    .o(al_3ca44efd[22]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_5880740 (
    .a(al_f2330f79[23]),
    .b(al_df7b4407),
    .o(al_3ca44efd[23]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_18cd1e72 (
    .a(al_f2330f79[24]),
    .b(al_df7b4407),
    .o(al_3ca44efd[24]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_6ab2d088 (
    .a(al_f2330f79[25]),
    .b(al_df7b4407),
    .o(al_3ca44efd[25]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_5ebdcff2 (
    .a(al_f2330f79[26]),
    .b(al_df7b4407),
    .o(al_3ca44efd[26]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_e54aec11 (
    .a(al_f2330f79[27]),
    .b(al_df7b4407),
    .o(al_3ca44efd[27]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_22f99786 (
    .a(al_f2330f79[28]),
    .b(al_df7b4407),
    .o(al_3ca44efd[28]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_9d999b0a (
    .a(al_f2330f79[29]),
    .b(al_df7b4407),
    .o(al_3ca44efd[29]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_e08fa253 (
    .a(al_f2330f79[2]),
    .b(al_df7b4407),
    .o(al_3ca44efd[2]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_d64d3ae (
    .a(al_f2330f79[30]),
    .b(al_df7b4407),
    .o(al_3ca44efd[30]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_dc9b560b (
    .a(al_f2330f79[31]),
    .b(al_df7b4407),
    .o(al_3ca44efd[31]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_3502b7c9 (
    .a(al_f2330f79[3]),
    .b(al_df7b4407),
    .o(al_3ca44efd[3]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_47b9c0f2 (
    .a(al_f2330f79[4]),
    .b(al_df7b4407),
    .o(al_3ca44efd[4]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_6f291644 (
    .a(al_f2330f79[5]),
    .b(al_df7b4407),
    .o(al_3ca44efd[5]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_e0c559b0 (
    .a(al_f2330f79[6]),
    .b(al_df7b4407),
    .o(al_3ca44efd[6]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_e8b5de3d (
    .a(al_f2330f79[7]),
    .b(al_df7b4407),
    .o(al_3ca44efd[7]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_3fbfad47 (
    .a(al_f2330f79[8]),
    .b(al_df7b4407),
    .o(al_3ca44efd[8]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_7b1a06e9 (
    .a(al_f2330f79[9]),
    .b(al_df7b4407),
    .o(al_3ca44efd[9]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_f980b0d9 (
    .a(al_9d63e9cd),
    .b(al_6ec8afa5),
    .o(al_1a1af7e4));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_47849044 (
    .a(al_6a0e908c),
    .b(al_5e60a110),
    .c(al_6ec8afa5),
    .o(al_119831c0));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    al_1ba2d6b8 (
    .a(al_c795a432),
    .b(al_a8151162),
    .c(al_7d2c853e),
    .o(al_66ffb9));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9139c1d1 (
    .a(al_a7b01c14[2]),
    .b(al_c46301d),
    .o(al_a25a6119));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_4fed55ba (
    .a(al_1a1af7e4),
    .b(al_119831c0),
    .c(al_6a6f79fc),
    .o(al_c83b3308));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*~(~C*B*A)))*~(D)+~F*(~E*~(~C*B*A))*~(D)+~(~F)*(~E*~(~C*B*A))*D+~F*(~E*~(~C*B*A))*D)"),
    .INIT(64'hffff08ffff000800))
    al_a0365310 (
    .a(al_a25a6119),
    .b(al_c83b3308),
    .c(al_66ffb9),
    .d(iBusAhb_HREADY),
    .e(al_48d2ef94),
    .f(al_a4f21dd7),
    .o(al_589bdcdb));
  AL_DFF_X al_7b2fce8 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_589bdcdb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a4f21dd7));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f3b7cd1c (
    .a(al_a0e6869c[13]),
    .b(al_7b59c46e[0]),
    .c(al_b70cb9be[0]),
    .o(al_94f1da4c[0]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_3c981bd2 (
    .a(al_94f1da4c[0]),
    .b(al_a167c8cf),
    .o(al_f3b8f942[0]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_e5f10ec6 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[10]),
    .d(al_b70cb9be[10]),
    .o(al_f3b8f942[10]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_8b607d55 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[11]),
    .d(al_b70cb9be[11]),
    .o(al_f3b8f942[11]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_db2e28b8 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[12]),
    .d(al_b70cb9be[12]),
    .o(al_f3b8f942[12]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_895e2618 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[13]),
    .d(al_b70cb9be[13]),
    .o(al_f3b8f942[13]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_20d6c2b9 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[14]),
    .d(al_b70cb9be[14]),
    .o(al_f3b8f942[14]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_9fc8241a (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[15]),
    .d(al_b70cb9be[15]),
    .o(al_f3b8f942[15]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_338d06f4 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[16]),
    .d(al_b70cb9be[16]),
    .o(al_f3b8f942[16]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_c0da8438 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[17]),
    .d(al_b70cb9be[17]),
    .o(al_f3b8f942[17]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_cec9f287 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[18]),
    .d(al_b70cb9be[18]),
    .o(al_f3b8f942[18]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_4bcf1cf3 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[19]),
    .d(al_b70cb9be[19]),
    .o(al_f3b8f942[19]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_a01c8964 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[1]),
    .d(al_b70cb9be[1]),
    .o(al_f3b8f942[1]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_f1c5e804 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[20]),
    .d(al_b70cb9be[20]),
    .o(al_f3b8f942[20]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_5d779e4d (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[21]),
    .d(al_b70cb9be[21]),
    .o(al_f3b8f942[21]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_4651d851 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[22]),
    .d(al_b70cb9be[22]),
    .o(al_f3b8f942[22]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_d4caa0df (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[23]),
    .d(al_b70cb9be[23]),
    .o(al_f3b8f942[23]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_9b90af8b (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[24]),
    .d(al_b70cb9be[24]),
    .o(al_f3b8f942[24]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_f70b1506 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[25]),
    .d(al_b70cb9be[25]),
    .o(al_f3b8f942[25]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_ff220796 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[26]),
    .d(al_b70cb9be[26]),
    .o(al_f3b8f942[26]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_b0e62c1d (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[27]),
    .d(al_b70cb9be[27]),
    .o(al_f3b8f942[27]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_2f68d13f (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[28]),
    .d(al_b70cb9be[28]),
    .o(al_f3b8f942[28]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_603b7847 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[29]),
    .d(al_b70cb9be[29]),
    .o(al_f3b8f942[29]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_43c2e2f3 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[2]),
    .d(al_b70cb9be[2]),
    .o(al_f3b8f942[2]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_eb68891c (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[30]),
    .d(al_b70cb9be[30]),
    .o(al_f3b8f942[30]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_45b4b047 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[31]),
    .d(al_b70cb9be[31]),
    .o(al_f3b8f942[31]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_abdad7f4 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[3]),
    .d(al_b70cb9be[3]),
    .o(al_f3b8f942[3]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_e3f2905a (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[4]),
    .d(al_b70cb9be[4]),
    .o(al_f3b8f942[4]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_a2daad4a (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[5]),
    .d(al_b70cb9be[5]),
    .o(al_f3b8f942[5]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_ebc65f86 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[6]),
    .d(al_b70cb9be[6]),
    .o(al_f3b8f942[6]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_5bc841b9 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[7]),
    .d(al_b70cb9be[7]),
    .o(al_f3b8f942[7]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_7eff91d1 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[8]),
    .d(al_b70cb9be[8]),
    .o(al_f3b8f942[8]));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h596a))
    al_24775cc0 (
    .a(al_a167c8cf),
    .b(al_a0e6869c[13]),
    .c(al_7b59c46e[9]),
    .d(al_b70cb9be[9]),
    .o(al_f3b8f942[9]));
  AL_DFF_X al_6b67c5da (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_4fdb397d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b8fe1a1f));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*A))*~(B)+C*(D*A)*~(B)+~(C)*(D*A)*B+C*(D*A)*B)"),
    .INIT(16'hb830))
    al_bf468ffa (
    .a(al_1a09507b),
    .b(dBusAhb_HREADY_IN),
    .c(al_b8fe1a1f),
    .d(dBusAhb_HWRITE),
    .o(al_4fdb397d));
  AL_DFF_X al_1e98c95a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d4a46bf1));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_c100b811 (
    .a(1'b0),
    .o({al_2672f5b2,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_486b583c (
    .a(al_a16ef20a[1]),
    .b(al_1d7074bf),
    .c(al_2672f5b2),
    .o({al_82ca9a92,al_e79b3dfa}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_183bdf14 (
    .a(al_a16ef20a[2]),
    .b(al_4cc97ac1),
    .c(al_82ca9a92),
    .o({al_879c97c5,al_ca581e6c}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f2646b7 (
    .a(al_a16ef20a[3]),
    .b(al_de666865),
    .c(al_879c97c5),
    .o({al_837e8da8,al_428b50b6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_53346e5a (
    .a(al_a16ef20a[4]),
    .b(al_a40c439),
    .c(al_837e8da8),
    .o({al_9c95e435,al_a3f3ee06}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_48a43b42 (
    .a(al_a16ef20a[5]),
    .b(al_85a2bdb0[25]),
    .c(al_9c95e435),
    .o({al_542d1ba4,al_263322e4}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e69a150 (
    .a(al_a16ef20a[6]),
    .b(al_85a2bdb0[26]),
    .c(al_542d1ba4),
    .o({al_f4e939bc,al_63bbd3a2}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5d7c35e2 (
    .a(al_a16ef20a[7]),
    .b(al_85a2bdb0[27]),
    .c(al_f4e939bc),
    .o({al_26903ef3,al_6ab73d4d}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_984f52c8 (
    .a(al_a16ef20a[8]),
    .b(al_85a2bdb0[28]),
    .c(al_26903ef3),
    .o({al_82a77528,al_fd8d8e0c}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_49264961 (
    .a(al_a16ef20a[9]),
    .b(al_85a2bdb0[29]),
    .c(al_82a77528),
    .o({al_5b477973,al_a89113a9}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d02ac232 (
    .a(al_a16ef20a[10]),
    .b(al_85a2bdb0[30]),
    .c(al_5b477973),
    .o({al_12fa803d,al_8d9bdfff}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9fceb363 (
    .a(al_a16ef20a[11]),
    .b(al_1405651f),
    .c(al_12fa803d),
    .o({al_6426fa0c,al_70f172be}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_53ef7dab (
    .a(al_a16ef20a[12]),
    .b(al_383f9835),
    .c(al_6426fa0c),
    .o({al_8b1fccb,al_c89d1229}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b0a7c58 (
    .a(al_a16ef20a[13]),
    .b(al_420d5318),
    .c(al_8b1fccb),
    .o({al_4e576557,al_2d354b}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9b508627 (
    .a(al_a16ef20a[14]),
    .b(al_2cce4860),
    .c(al_4e576557),
    .o({al_6c384295,al_2fb7633}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_88461592 (
    .a(al_a16ef20a[15]),
    .b(al_96c3cafb),
    .c(al_6c384295),
    .o({al_63a3bec2,al_5b3ba944}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_12120cb0 (
    .a(al_a16ef20a[16]),
    .b(al_bcf22cd5),
    .c(al_63a3bec2),
    .o({al_4a1a4a4,al_f5f3edb6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f380056f (
    .a(al_a16ef20a[17]),
    .b(al_4bfb7d3a),
    .c(al_4a1a4a4),
    .o({al_7f54ca49,al_d0702be9}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7d725d5d (
    .a(al_a16ef20a[18]),
    .b(al_cc14dad7),
    .c(al_7f54ca49),
    .o({al_16541a17,al_2eb5050b}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_213b3486 (
    .a(al_a16ef20a[19]),
    .b(al_8c22c3eb),
    .c(al_16541a17),
    .o({al_2bfbeb6,al_89a93b84}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cbf55361 (
    .a(al_a16ef20a[20]),
    .b(al_85a2bdb0[31]),
    .c(al_2bfbeb6),
    .o({al_1f8435f6,al_82b168eb}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bc64eb0b (
    .a(al_a16ef20a[21]),
    .b(al_85a2bdb0[31]),
    .c(al_1f8435f6),
    .o({al_24d740cb,al_e2259475}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a09aa8ef (
    .a(al_a16ef20a[22]),
    .b(al_85a2bdb0[31]),
    .c(al_24d740cb),
    .o({al_f2f80319,al_6758eae2}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5b219f52 (
    .a(al_a16ef20a[23]),
    .b(al_85a2bdb0[31]),
    .c(al_f2f80319),
    .o({al_80daf3e,al_f814979a}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_57d66a05 (
    .a(al_a16ef20a[24]),
    .b(al_85a2bdb0[31]),
    .c(al_80daf3e),
    .o({al_f50ab810,al_5ca98598}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3853e547 (
    .a(al_a16ef20a[25]),
    .b(al_85a2bdb0[31]),
    .c(al_f50ab810),
    .o({al_3d0077da,al_267d2aa}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_503efa84 (
    .a(al_a16ef20a[26]),
    .b(al_85a2bdb0[31]),
    .c(al_3d0077da),
    .o({al_73502252,al_debfa536}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f7c984a0 (
    .a(al_a16ef20a[27]),
    .b(al_85a2bdb0[31]),
    .c(al_73502252),
    .o({al_df3a7245,al_f19f190e}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6494be3 (
    .a(al_a16ef20a[28]),
    .b(al_85a2bdb0[31]),
    .c(al_df3a7245),
    .o({al_829d1309,al_9852e0df}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_40a54fe2 (
    .a(al_a16ef20a[29]),
    .b(al_85a2bdb0[31]),
    .c(al_829d1309),
    .o({al_966d08ce,al_ecd761fc}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ea6b3a54 (
    .a(al_a16ef20a[30]),
    .b(al_85a2bdb0[31]),
    .c(al_966d08ce),
    .o({al_d8039a59,al_c64cf9f6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_24c73c37 (
    .a(al_a16ef20a[31]),
    .b(al_85a2bdb0[31]),
    .c(al_d8039a59),
    .o({open_n15,al_5e07bd5e}));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_f1d1cda4 (
    .a(al_3d2fbc2e[33]),
    .b(al_9edb1d1e[33]),
    .c(1'b0),
    .o(al_8f26ae38[33]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_4704d6be (
    .a(al_ccb50b3a[16]),
    .b(al_3d2fbc2e[0]),
    .c(al_9edb1d1e[0]),
    .o(al_8b049eb2[1]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_17d3858d (
    .a(al_ccb50b3a[17]),
    .b(al_3d2fbc2e[1]),
    .c(al_9edb1d1e[1]),
    .o(al_8b049eb2[2]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_1c383563 (
    .a(al_ccb50b3a[18]),
    .b(al_3d2fbc2e[2]),
    .c(al_9edb1d1e[2]),
    .o(al_8b049eb2[3]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_92e2a3b (
    .a(al_ccb50b3a[19]),
    .b(al_3d2fbc2e[3]),
    .c(al_9edb1d1e[3]),
    .o(al_8b049eb2[4]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_fc59cf0b (
    .a(al_ccb50b3a[20]),
    .b(al_3d2fbc2e[4]),
    .c(al_9edb1d1e[4]),
    .o(al_8b049eb2[5]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_636c4ce7 (
    .a(al_ccb50b3a[21]),
    .b(al_3d2fbc2e[5]),
    .c(al_9edb1d1e[5]),
    .o(al_8b049eb2[6]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_ecc7a994 (
    .a(al_ccb50b3a[22]),
    .b(al_3d2fbc2e[6]),
    .c(al_9edb1d1e[6]),
    .o(al_8b049eb2[7]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_73c0cdba (
    .a(al_ccb50b3a[23]),
    .b(al_3d2fbc2e[7]),
    .c(al_9edb1d1e[7]),
    .o(al_8b049eb2[8]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_9ecb11d (
    .a(al_ccb50b3a[24]),
    .b(al_3d2fbc2e[8]),
    .c(al_9edb1d1e[8]),
    .o(al_8b049eb2[9]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_9c75cb8b (
    .a(al_ccb50b3a[25]),
    .b(al_3d2fbc2e[9]),
    .c(al_9edb1d1e[9]),
    .o(al_8b049eb2[10]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_9815fcc2 (
    .a(al_ccb50b3a[26]),
    .b(al_3d2fbc2e[10]),
    .c(al_9edb1d1e[10]),
    .o(al_8b049eb2[11]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_50d95bde (
    .a(al_ccb50b3a[27]),
    .b(al_3d2fbc2e[11]),
    .c(al_9edb1d1e[11]),
    .o(al_8b049eb2[12]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_b32f5555 (
    .a(al_ccb50b3a[28]),
    .b(al_3d2fbc2e[12]),
    .c(al_9edb1d1e[12]),
    .o(al_8b049eb2[13]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_84eab8de (
    .a(al_ccb50b3a[29]),
    .b(al_3d2fbc2e[13]),
    .c(al_9edb1d1e[13]),
    .o(al_8b049eb2[14]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_e6fe02f7 (
    .a(al_ccb50b3a[30]),
    .b(al_3d2fbc2e[14]),
    .c(al_9edb1d1e[14]),
    .o(al_8b049eb2[15]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_cc558593 (
    .a(al_ccb50b3a[31]),
    .b(al_3d2fbc2e[15]),
    .c(al_9edb1d1e[15]),
    .o(al_8b049eb2[16]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_8bfc92a9 (
    .a(al_3d2fbc2e[16]),
    .b(al_9edb1d1e[16]),
    .c(1'b0),
    .o(al_8b049eb2[17]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_e1755951 (
    .a(al_3d2fbc2e[17]),
    .b(al_9edb1d1e[17]),
    .c(1'b0),
    .o(al_8b049eb2[18]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_e8eb52d4 (
    .a(al_3d2fbc2e[18]),
    .b(al_9edb1d1e[18]),
    .c(1'b0),
    .o(al_8b049eb2[19]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_743f771b (
    .a(al_3d2fbc2e[19]),
    .b(al_9edb1d1e[19]),
    .c(1'b0),
    .o(al_8b049eb2[20]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_970a3d38 (
    .a(al_3d2fbc2e[20]),
    .b(al_9edb1d1e[20]),
    .c(1'b0),
    .o(al_8b049eb2[21]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_e6593dd7 (
    .a(al_3d2fbc2e[21]),
    .b(al_9edb1d1e[21]),
    .c(1'b0),
    .o(al_8b049eb2[22]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_dc2cd6c6 (
    .a(al_3d2fbc2e[22]),
    .b(al_9edb1d1e[22]),
    .c(1'b0),
    .o(al_8b049eb2[23]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_6a52558c (
    .a(al_3d2fbc2e[23]),
    .b(al_9edb1d1e[23]),
    .c(1'b0),
    .o(al_8b049eb2[24]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_eee8c5af (
    .a(al_3d2fbc2e[24]),
    .b(al_9edb1d1e[24]),
    .c(1'b0),
    .o(al_8b049eb2[25]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_44502d0a (
    .a(al_3d2fbc2e[25]),
    .b(al_9edb1d1e[25]),
    .c(1'b0),
    .o(al_8b049eb2[26]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_d433531 (
    .a(al_3d2fbc2e[26]),
    .b(al_9edb1d1e[26]),
    .c(1'b0),
    .o(al_8b049eb2[27]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_2fdfb687 (
    .a(al_3d2fbc2e[27]),
    .b(al_9edb1d1e[27]),
    .c(1'b0),
    .o(al_8b049eb2[28]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_38d9a6a5 (
    .a(al_3d2fbc2e[28]),
    .b(al_9edb1d1e[28]),
    .c(1'b0),
    .o(al_8b049eb2[29]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_76d9a6fd (
    .a(al_3d2fbc2e[29]),
    .b(al_9edb1d1e[29]),
    .c(1'b0),
    .o(al_8b049eb2[30]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_f586f0a0 (
    .a(al_3d2fbc2e[30]),
    .b(al_9edb1d1e[30]),
    .c(1'b0),
    .o(al_8b049eb2[31]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_ac9e9120 (
    .a(al_3d2fbc2e[31]),
    .b(al_9edb1d1e[31]),
    .c(1'b0),
    .o(al_8b049eb2[32]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_17681b6 (
    .a(al_3d2fbc2e[32]),
    .b(al_9edb1d1e[32]),
    .c(1'b0),
    .o(al_8b049eb2[33]));
  AL_MAP_LUT3 #(
    .EQN("((A+B)*(A+C)*(B+C))"),
    .INIT(8'b11101000))
    al_8c2c0798 (
    .a(al_3d2fbc2e[33]),
    .b(al_9edb1d1e[33]),
    .c(1'b0),
    .o(al_8b049eb2[34]));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_5ca37f17 (
    .a(1'b0),
    .o({al_468d3b3e[1],open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dc863ec5 (
    .a(al_8f26ae38[1]),
    .b(al_8b049eb2[1]),
    .c(al_468d3b3e[1]),
    .o({al_468d3b3e[2],al_8dd2d746[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7abb49c4 (
    .a(al_8f26ae38[2]),
    .b(al_8b049eb2[2]),
    .c(al_468d3b3e[2]),
    .o({al_468d3b3e[3],al_8dd2d746[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ed01b0c7 (
    .a(al_8f26ae38[3]),
    .b(al_8b049eb2[3]),
    .c(al_468d3b3e[3]),
    .o({al_468d3b3e[4],al_8dd2d746[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5a27bd55 (
    .a(al_8f26ae38[4]),
    .b(al_8b049eb2[4]),
    .c(al_468d3b3e[4]),
    .o({al_468d3b3e[5],al_8dd2d746[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_52521482 (
    .a(al_8f26ae38[5]),
    .b(al_8b049eb2[5]),
    .c(al_468d3b3e[5]),
    .o({al_468d3b3e[6],al_8dd2d746[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f70613b1 (
    .a(al_8f26ae38[6]),
    .b(al_8b049eb2[6]),
    .c(al_468d3b3e[6]),
    .o({al_468d3b3e[7],al_8dd2d746[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6b2b7f17 (
    .a(al_8f26ae38[7]),
    .b(al_8b049eb2[7]),
    .c(al_468d3b3e[7]),
    .o({al_468d3b3e[8],al_8dd2d746[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e25d9f0e (
    .a(al_8f26ae38[8]),
    .b(al_8b049eb2[8]),
    .c(al_468d3b3e[8]),
    .o({al_468d3b3e[9],al_8dd2d746[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f724ebd (
    .a(al_8f26ae38[9]),
    .b(al_8b049eb2[9]),
    .c(al_468d3b3e[9]),
    .o({al_468d3b3e[10],al_8dd2d746[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8869da8 (
    .a(al_8f26ae38[10]),
    .b(al_8b049eb2[10]),
    .c(al_468d3b3e[10]),
    .o({al_468d3b3e[11],al_8dd2d746[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d4e5a95b (
    .a(al_8f26ae38[11]),
    .b(al_8b049eb2[11]),
    .c(al_468d3b3e[11]),
    .o({al_468d3b3e[12],al_8dd2d746[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3811b071 (
    .a(al_8f26ae38[12]),
    .b(al_8b049eb2[12]),
    .c(al_468d3b3e[12]),
    .o({al_468d3b3e[13],al_8dd2d746[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_76ebecaa (
    .a(al_8f26ae38[13]),
    .b(al_8b049eb2[13]),
    .c(al_468d3b3e[13]),
    .o({al_468d3b3e[14],al_8dd2d746[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_db80a1f8 (
    .a(al_8f26ae38[14]),
    .b(al_8b049eb2[14]),
    .c(al_468d3b3e[14]),
    .o({al_468d3b3e[15],al_8dd2d746[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ef48217e (
    .a(al_8f26ae38[15]),
    .b(al_8b049eb2[15]),
    .c(al_468d3b3e[15]),
    .o({al_468d3b3e[16],al_8dd2d746[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b5aedd3e (
    .a(al_8f26ae38[16]),
    .b(al_8b049eb2[16]),
    .c(al_468d3b3e[16]),
    .o({al_468d3b3e[17],al_8dd2d746[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_933d5579 (
    .a(al_8f26ae38[17]),
    .b(al_8b049eb2[17]),
    .c(al_468d3b3e[17]),
    .o({al_468d3b3e[18],al_8dd2d746[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3c3748a3 (
    .a(al_8f26ae38[18]),
    .b(al_8b049eb2[18]),
    .c(al_468d3b3e[18]),
    .o({al_468d3b3e[19],al_8dd2d746[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ea87a456 (
    .a(al_8f26ae38[19]),
    .b(al_8b049eb2[19]),
    .c(al_468d3b3e[19]),
    .o({al_468d3b3e[20],al_8dd2d746[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3ee313fa (
    .a(al_8f26ae38[20]),
    .b(al_8b049eb2[20]),
    .c(al_468d3b3e[20]),
    .o({al_468d3b3e[21],al_8dd2d746[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_15030cb7 (
    .a(al_8f26ae38[21]),
    .b(al_8b049eb2[21]),
    .c(al_468d3b3e[21]),
    .o({al_468d3b3e[22],al_8dd2d746[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_18c877b0 (
    .a(al_8f26ae38[22]),
    .b(al_8b049eb2[22]),
    .c(al_468d3b3e[22]),
    .o({al_468d3b3e[23],al_8dd2d746[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cc75118c (
    .a(al_8f26ae38[23]),
    .b(al_8b049eb2[23]),
    .c(al_468d3b3e[23]),
    .o({al_468d3b3e[24],al_8dd2d746[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_794e6bec (
    .a(al_8f26ae38[24]),
    .b(al_8b049eb2[24]),
    .c(al_468d3b3e[24]),
    .o({al_468d3b3e[25],al_8dd2d746[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9f100eee (
    .a(al_8f26ae38[25]),
    .b(al_8b049eb2[25]),
    .c(al_468d3b3e[25]),
    .o({al_468d3b3e[26],al_8dd2d746[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f5e02581 (
    .a(al_8f26ae38[26]),
    .b(al_8b049eb2[26]),
    .c(al_468d3b3e[26]),
    .o({al_468d3b3e[27],al_8dd2d746[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cb01ae78 (
    .a(al_8f26ae38[27]),
    .b(al_8b049eb2[27]),
    .c(al_468d3b3e[27]),
    .o({al_468d3b3e[28],al_8dd2d746[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8f9cf891 (
    .a(al_8f26ae38[28]),
    .b(al_8b049eb2[28]),
    .c(al_468d3b3e[28]),
    .o({al_468d3b3e[29],al_8dd2d746[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8d0f9c86 (
    .a(al_8f26ae38[29]),
    .b(al_8b049eb2[29]),
    .c(al_468d3b3e[29]),
    .o({al_468d3b3e[30],al_8dd2d746[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e4a5be67 (
    .a(al_8f26ae38[30]),
    .b(al_8b049eb2[30]),
    .c(al_468d3b3e[30]),
    .o({al_468d3b3e[31],al_8dd2d746[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_279b5688 (
    .a(al_8f26ae38[31]),
    .b(al_8b049eb2[31]),
    .c(al_468d3b3e[31]),
    .o({al_468d3b3e[32],al_8dd2d746[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7c8e6a79 (
    .a(al_8f26ae38[32]),
    .b(al_8b049eb2[32]),
    .c(al_468d3b3e[32]),
    .o({al_468d3b3e[33],al_8dd2d746[32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_872aa286 (
    .a(al_8f26ae38[33]),
    .b(al_8b049eb2[33]),
    .c(al_468d3b3e[33]),
    .o({al_468d3b3e[34],al_8dd2d746[33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b41554fd (
    .a(al_8f26ae38[33]),
    .b(al_8b049eb2[34]),
    .c(al_468d3b3e[34]),
    .o({al_468d3b3e[35],al_8dd2d746[34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_809da70a (
    .a(al_8f26ae38[33]),
    .b(al_8b049eb2[34]),
    .c(al_468d3b3e[35]),
    .o({open_n19,al_8dd2d746[35]}));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_6f31f2fd (
    .a(al_ccb50b3a[16]),
    .b(al_3d2fbc2e[0]),
    .c(al_9edb1d1e[0]),
    .o(al_8dd2d746[0]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_5ac58c7 (
    .a(al_ccb50b3a[17]),
    .b(al_3d2fbc2e[1]),
    .c(al_9edb1d1e[1]),
    .o(al_8f26ae38[1]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_d2c61aea (
    .a(al_ccb50b3a[18]),
    .b(al_3d2fbc2e[2]),
    .c(al_9edb1d1e[2]),
    .o(al_8f26ae38[2]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_b941fe7b (
    .a(al_ccb50b3a[19]),
    .b(al_3d2fbc2e[3]),
    .c(al_9edb1d1e[3]),
    .o(al_8f26ae38[3]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_193b185c (
    .a(al_ccb50b3a[20]),
    .b(al_3d2fbc2e[4]),
    .c(al_9edb1d1e[4]),
    .o(al_8f26ae38[4]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_b2f5017a (
    .a(al_ccb50b3a[21]),
    .b(al_3d2fbc2e[5]),
    .c(al_9edb1d1e[5]),
    .o(al_8f26ae38[5]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_7c0a44e2 (
    .a(al_ccb50b3a[22]),
    .b(al_3d2fbc2e[6]),
    .c(al_9edb1d1e[6]),
    .o(al_8f26ae38[6]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_ff3c82e7 (
    .a(al_ccb50b3a[23]),
    .b(al_3d2fbc2e[7]),
    .c(al_9edb1d1e[7]),
    .o(al_8f26ae38[7]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_574508b (
    .a(al_ccb50b3a[24]),
    .b(al_3d2fbc2e[8]),
    .c(al_9edb1d1e[8]),
    .o(al_8f26ae38[8]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_954ca94f (
    .a(al_ccb50b3a[25]),
    .b(al_3d2fbc2e[9]),
    .c(al_9edb1d1e[9]),
    .o(al_8f26ae38[9]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_2a1864cb (
    .a(al_ccb50b3a[26]),
    .b(al_3d2fbc2e[10]),
    .c(al_9edb1d1e[10]),
    .o(al_8f26ae38[10]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_59251cb3 (
    .a(al_ccb50b3a[27]),
    .b(al_3d2fbc2e[11]),
    .c(al_9edb1d1e[11]),
    .o(al_8f26ae38[11]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_ec034541 (
    .a(al_ccb50b3a[28]),
    .b(al_3d2fbc2e[12]),
    .c(al_9edb1d1e[12]),
    .o(al_8f26ae38[12]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_f1e23351 (
    .a(al_ccb50b3a[29]),
    .b(al_3d2fbc2e[13]),
    .c(al_9edb1d1e[13]),
    .o(al_8f26ae38[13]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_41904c6c (
    .a(al_ccb50b3a[30]),
    .b(al_3d2fbc2e[14]),
    .c(al_9edb1d1e[14]),
    .o(al_8f26ae38[14]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_a07a3c1 (
    .a(al_ccb50b3a[31]),
    .b(al_3d2fbc2e[15]),
    .c(al_9edb1d1e[15]),
    .o(al_8f26ae38[15]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_d7dab6dc (
    .a(al_3d2fbc2e[16]),
    .b(al_9edb1d1e[16]),
    .c(1'b0),
    .o(al_8f26ae38[16]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_836df61c (
    .a(al_3d2fbc2e[17]),
    .b(al_9edb1d1e[17]),
    .c(1'b0),
    .o(al_8f26ae38[17]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_2a30a6f6 (
    .a(al_3d2fbc2e[18]),
    .b(al_9edb1d1e[18]),
    .c(1'b0),
    .o(al_8f26ae38[18]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_5f51d72f (
    .a(al_3d2fbc2e[19]),
    .b(al_9edb1d1e[19]),
    .c(1'b0),
    .o(al_8f26ae38[19]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_1cf0af06 (
    .a(al_3d2fbc2e[20]),
    .b(al_9edb1d1e[20]),
    .c(1'b0),
    .o(al_8f26ae38[20]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_2e122ad4 (
    .a(al_3d2fbc2e[21]),
    .b(al_9edb1d1e[21]),
    .c(1'b0),
    .o(al_8f26ae38[21]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_eb82939a (
    .a(al_3d2fbc2e[22]),
    .b(al_9edb1d1e[22]),
    .c(1'b0),
    .o(al_8f26ae38[22]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_5bb2089a (
    .a(al_3d2fbc2e[23]),
    .b(al_9edb1d1e[23]),
    .c(1'b0),
    .o(al_8f26ae38[23]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_589531e (
    .a(al_3d2fbc2e[24]),
    .b(al_9edb1d1e[24]),
    .c(1'b0),
    .o(al_8f26ae38[24]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_25ee8f1f (
    .a(al_3d2fbc2e[25]),
    .b(al_9edb1d1e[25]),
    .c(1'b0),
    .o(al_8f26ae38[25]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_8d1ce725 (
    .a(al_3d2fbc2e[26]),
    .b(al_9edb1d1e[26]),
    .c(1'b0),
    .o(al_8f26ae38[26]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_371f485 (
    .a(al_3d2fbc2e[27]),
    .b(al_9edb1d1e[27]),
    .c(1'b0),
    .o(al_8f26ae38[27]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_9adb0082 (
    .a(al_3d2fbc2e[28]),
    .b(al_9edb1d1e[28]),
    .c(1'b0),
    .o(al_8f26ae38[28]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_47839a83 (
    .a(al_3d2fbc2e[29]),
    .b(al_9edb1d1e[29]),
    .c(1'b0),
    .o(al_8f26ae38[29]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_8f490ae3 (
    .a(al_3d2fbc2e[30]),
    .b(al_9edb1d1e[30]),
    .c(1'b0),
    .o(al_8f26ae38[30]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_65822a64 (
    .a(al_3d2fbc2e[31]),
    .b(al_9edb1d1e[31]),
    .c(1'b0),
    .o(al_8f26ae38[31]));
  AL_MAP_LUT3 #(
    .EQN("(A@B@C)"),
    .INIT(8'b10010110))
    al_a8d7e08a (
    .a(al_3d2fbc2e[32]),
    .b(al_9edb1d1e[32]),
    .c(1'b0),
    .o(al_8f26ae38[32]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_f8d64848 (
    .a(al_6faa66d6),
    .b(al_85a2bdb0[18]),
    .c(al_85a2bdb0[19]),
    .d(al_e03b3126[10]),
    .e(al_e03b3126[11]),
    .o(al_a62203af));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc0c3c1438087c547))
    al_67c576e0 (
    .a(al_85a2bdb0[4]),
    .b(al_85a2bdb0[5]),
    .c(al_85a2bdb0[6]),
    .d(al_85a2bdb0[12]),
    .e(al_85a2bdb0[13]),
    .f(al_85a2bdb0[14]),
    .o(al_c6d62120));
  AL_MAP_LUT6 #(
    .EQN("(F*~(~C*~(D@B)*~(E*A)))"),
    .INIT(64'hfbfef3fc00000000))
    al_6a03ae98 (
    .a(al_85a2bdb0[5]),
    .b(al_85a2bdb0[12]),
    .c(al_85a2bdb0[13]),
    .d(al_85a2bdb0[14]),
    .e(al_85a2bdb0[25]),
    .f(al_85a2bdb0[30]),
    .o(al_2e313516));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_abeb0aa5 (
    .a(al_85a2bdb0[4]),
    .b(al_85a2bdb0[6]),
    .c(al_85a2bdb0[26]),
    .d(al_85a2bdb0[27]),
    .e(al_85a2bdb0[28]),
    .f(al_85a2bdb0[29]),
    .o(al_2f2822d8));
  AL_MAP_LUT6 #(
    .EQN("(~E*~D*~(~A*~(~F*C*~B)))"),
    .INIT(64'h000000aa000000ba))
    al_ddfb48ff (
    .a(al_c6d62120),
    .b(al_2e313516),
    .c(al_2f2822d8),
    .d(al_85a2bdb0[2]),
    .e(al_85a2bdb0[3]),
    .f(al_85a2bdb0[31]),
    .o(al_99aa8cdf));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf7ffdfcff7ffdfdf))
    al_cfa53f35 (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[3]),
    .c(al_85a2bdb0[4]),
    .d(al_85a2bdb0[5]),
    .e(al_85a2bdb0[6]),
    .f(al_85a2bdb0[13]),
    .o(al_2a7e21ae));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*~A))"),
    .INIT(16'hb000))
    al_1aa245d7 (
    .a(al_99aa8cdf),
    .b(al_2a7e21ae),
    .c(al_85a2bdb0[0]),
    .d(al_85a2bdb0[1]),
    .o(al_26f3954d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_58a5c2c1 (
    .a(al_85a2bdb0[0]),
    .b(al_85a2bdb0[1]),
    .c(al_85a2bdb0[26]),
    .d(al_85a2bdb0[27]),
    .e(al_85a2bdb0[30]),
    .f(al_85a2bdb0[31]),
    .o(al_e4d5d147));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_c4fe6021 (
    .a(al_e4d5d147),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[14]),
    .d(al_85a2bdb0[19]),
    .e(al_85a2bdb0[23]),
    .o(al_c0f96426));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~D*~C*B*A)"),
    .INIT(64'h0008000000000000))
    al_9fff18ba (
    .a(al_c0f96426),
    .b(al_1a551855),
    .c(al_85a2bdb0[2]),
    .d(al_85a2bdb0[3]),
    .e(al_85a2bdb0[5]),
    .f(al_85a2bdb0[6]),
    .o(al_8b7c83a7));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_a5f2c435 (
    .a(al_85a2bdb0[15]),
    .b(al_85a2bdb0[16]),
    .c(al_85a2bdb0[17]),
    .d(al_85a2bdb0[18]),
    .e(al_85a2bdb0[24]),
    .f(al_85a2bdb0[25]),
    .o(al_95a8aeaf));
  AL_MAP_LUT6 #(
    .EQN("(A*(~(B)*~(C)*~(D)*~(E)*~(F)+B*~(C)*~(D)*~(E)*~(F)+~(B)*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+~(B)*C*~(D)*E*F))"),
    .INIT(64'h002000000820000a))
    al_4af2c75b (
    .a(al_95a8aeaf),
    .b(al_85a2bdb0[20]),
    .c(al_85a2bdb0[21]),
    .d(al_85a2bdb0[22]),
    .e(al_85a2bdb0[28]),
    .f(al_85a2bdb0[29]),
    .o(al_4be831c2));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_efbd7bd6 (
    .a(al_85a2bdb0[0]),
    .b(al_85a2bdb0[1]),
    .c(al_85a2bdb0[4]),
    .d(al_85a2bdb0[13]),
    .e(al_85a2bdb0[14]),
    .o(al_277cf2f2));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*C*~(D)*~(E)*~(F)+~(B)*~(C)*D*E*~(F)+B*~(C)*D*E*~(F)+B*C*~(D)*~(E)*F))"),
    .INIT(64'h000000800a000080))
    al_44daf7ec (
    .a(al_277cf2f2),
    .b(al_85a2bdb0[2]),
    .c(al_85a2bdb0[3]),
    .d(al_85a2bdb0[5]),
    .e(al_85a2bdb0[6]),
    .f(al_85a2bdb0[12]),
    .o(al_8ac7c093));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_2ac0581c (
    .a(al_f49992c3),
    .b(al_202f2c67[0]),
    .c(al_202f2c67[1]),
    .d(al_202f2c67[2]),
    .o(al_c76629d2));
  AL_MAP_LUT6 #(
    .EQN("(~D*A*((C*B)*~(E)*~(F)+(C*B)*E*~(F)+~((C*B))*E*F+(C*B)*E*F))"),
    .INIT(64'h00aa000000800080))
    al_447be5a9 (
    .a(al_c76629d2),
    .b(al_acd38e8e),
    .c(iBusAhb_HRESP),
    .d(al_c73c0ba3),
    .e(al_b86dd14b[0]),
    .f(al_d518b626),
    .o(al_a3a8b68d));
  AL_MAP_LUT6 #(
    .EQN("(~E*~(~F*~D*~A*~(C*B)))"),
    .INIT(64'h0000ffff0000ffea))
    al_cc19ab38 (
    .a(al_26f3954d),
    .b(al_8b7c83a7),
    .c(al_4be831c2),
    .d(al_8ac7c093),
    .e(al_a3a8b68d),
    .f(al_f6cd735f),
    .o(al_a8151162));
  AL_MAP_LUT6 #(
    .EQN("(~F*~(A*~(~E*~D*~C*~B)))"),
    .INIT(64'h0000000055555557))
    al_e3b7eaaa (
    .a(al_6715e869),
    .b(al_235de557),
    .c(al_9c55c5c3),
    .d(al_4cc0b8dd),
    .e(al_7610b7fc),
    .f(al_809b319),
    .o(al_11418f51));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_53d02d05 (
    .a(al_e9897485),
    .b(al_804ebeec),
    .c(al_d19b9f6b),
    .d(al_be8ea5e1),
    .o(al_f170970d));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_b3386279 (
    .a(al_523cde28),
    .b(al_b5f1afb5[0]),
    .c(al_b5f1afb5[1]),
    .o(al_c85db05d));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*B*A))"),
    .INIT(16'h070f))
    al_da65d95 (
    .a(al_11418f51),
    .b(al_f170970d),
    .c(al_c85db05d),
    .d(al_b211b12d),
    .o(al_a5849610));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    al_6b8b58e5 (
    .a(al_5e275e81),
    .b(al_cbdc72d2),
    .c(al_cd3d5e6f),
    .d(al_501dbbdf),
    .o(al_12227f77));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    al_29f291fa (
    .a(al_1d840c32),
    .b(al_12227f77),
    .c(al_a430e4d2),
    .d(al_ea2eaeb1),
    .o(al_c572d1c7));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    al_b5172d79 (
    .a(al_c91705db),
    .b(al_ea2eaeb1),
    .c(al_cd3d5e6f),
    .d(al_501dbbdf),
    .o(al_6a0e908c));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_b149f693 (
    .a(al_6a0e908c),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e379ebb5),
    .e(al_a2deaa78),
    .o(al_c795a432));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    al_ab902b6a (
    .a(al_f6cd735f),
    .b(al_b567677b),
    .c(al_6893b11d),
    .d(al_69807e37),
    .o(al_c197c567));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_92149ac1 (
    .a(al_da9c21fb),
    .b(al_f6cd735f),
    .o(al_2c3e73df));
  AL_MAP_LUT6 #(
    .EQN("(D*~(~F*E*C*~B*~A))"),
    .INIT(64'hff00ff00ef00ff00))
    al_5084889f (
    .a(al_bec39e4d),
    .b(al_6ec8afa5),
    .c(al_c572d1c7),
    .d(dBusAhb_HREADY_IN),
    .e(al_b8fe1a1f),
    .f(dBusAhb_HWRITE),
    .o(al_291d5f8b));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~A*~(E*~D*~B)))"),
    .INIT(32'ha0b0a0a0))
    al_24564bf1 (
    .a(al_cbdc72d2),
    .b(al_bb6ca07d),
    .c(al_523cde28),
    .d(al_b5f1afb5[0]),
    .e(al_b5f1afb5[1]),
    .o(al_cdfe2d97));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*~(C*~(~E*~D)))"),
    .INIT(32'h02020222))
    al_5f368eb6 (
    .a(al_bb0cd305),
    .b(al_cdfe2d97),
    .c(al_b211b12d),
    .d(al_501dbbdf),
    .e(al_c0a7a5f),
    .o(al_71fb98b4));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E*D*~B*~A))"),
    .INIT(32'he0f0f0f0))
    al_eaa4c19a (
    .a(al_291d5f8b),
    .b(al_7bc36116),
    .c(al_71fb98b4),
    .d(al_32fedef4),
    .e(al_523cde28),
    .o(al_5a744f0f));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    al_da50cbe4 (
    .a(al_a5849610),
    .b(al_e379ebb5),
    .c(al_b469f7cc),
    .o(al_5e60a110));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    al_bc3cd9d5 (
    .a(al_de0f70d9),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[6]),
    .o(al_4f6deaed));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_5cf881d1 (
    .a(al_ebace85),
    .b(al_44595135),
    .c(al_523cde28),
    .o(al_3e5baa1a));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_801ee5ca (
    .a(al_cdace779),
    .b(al_24641d37),
    .c(al_501dbbdf),
    .o(al_5bcb7210));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    al_474dfe2e (
    .a(al_358f5bea),
    .b(al_df2df2f9),
    .c(al_4f6deaed),
    .d(al_3e5baa1a),
    .e(al_5bcb7210),
    .o(al_f66ced67));
  AL_MAP_LUT6 #(
    .EQN("(~(~D*~C)*~(~B*~(E*~(~F*~A))))"),
    .INIT(64'hfff0ccc0eee0ccc0))
    al_cca1c43f (
    .a(al_8bea08a7),
    .b(al_85a2bdb0[2]),
    .c(al_85a2bdb0[3]),
    .d(al_85a2bdb0[4]),
    .e(al_85a2bdb0[6]),
    .f(al_85a2bdb0[14]),
    .o(al_7167debf));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~(E*B)*~(D*A)))"),
    .INIT(32'h0e0c0a00))
    al_7c70fa06 (
    .a(al_a62203af),
    .b(al_a2426a1),
    .c(al_7167debf),
    .d(al_3e5baa1a),
    .e(al_5bcb7210),
    .o(al_ddfd7daa));
  AL_MAP_LUT6 #(
    .EQN("(~(~F*E*~D)*~(~C*B*A))"),
    .INIT(64'hf7f7f7f7f700f7f7))
    al_3856c54e (
    .a(al_523cde28),
    .b(al_b5f1afb5[0]),
    .c(al_b5f1afb5[1]),
    .d(al_5c72a609[0]),
    .e(al_5c72a609[1]),
    .f(al_5c72a609[2]),
    .o(al_134ffa88));
  AL_MAP_LUT6 #(
    .EQN("(~C*B*~A*~(~F*E*D))"),
    .INIT(64'h0404040400040404))
    al_ce22a18a (
    .a(al_c197c567),
    .b(al_134ffa88),
    .c(al_ea2eaeb1),
    .d(al_501dbbdf),
    .e(al_53188262[0]),
    .f(al_53188262[1]),
    .o(al_33a34bec));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(~B*~A)))"),
    .INIT(16'hf010))
    al_b9b53d40 (
    .a(al_f66ced67),
    .b(al_ddfd7daa),
    .c(al_33a34bec),
    .d(al_f6cd735f),
    .o(al_6f08d701));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_61ddd00b (
    .a(al_5a744f0f),
    .b(al_6f08d701),
    .o(al_a7b01c14[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_27d608f1 (
    .a(iBusAhb_HRDATA[0]),
    .b(al_b86dd14b[1]),
    .c(al_d518b626),
    .o(al_dc5d601));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cc208e4e (
    .a(iBusAhb_HRDATA[1]),
    .b(al_b86dd14b[2]),
    .c(al_d518b626),
    .o(al_39d0a986));
  AL_MAP_LUT6 #(
    .EQN("(E*D*A*~(~F*~(~C*~B)))"),
    .INIT(64'haa00000002000000))
    al_ffb020b0 (
    .a(al_5a744f0f),
    .b(al_f66ced67),
    .c(al_ddfd7daa),
    .d(al_33a34bec),
    .e(al_bd9d7d67),
    .f(al_f6cd735f),
    .o(al_1d3bfd2e));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_acad9416 (
    .a(al_cf18c1c6[16]),
    .b(al_cf18c1c6[17]),
    .o(al_d72f4570));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_e84764f6 (
    .a(al_dc5d601),
    .b(al_39d0a986),
    .o(al_fccc3291));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~C*~(~E*~D*~B)))"),
    .INIT(32'h50505051))
    al_3d0b2cce (
    .a(al_d72f4570),
    .b(al_fccc3291),
    .c(al_bccf82af),
    .d(al_9c16c2f5),
    .e(al_126b3afd[1]),
    .o(al_37a2cec8));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    al_648e5ef1 (
    .a(al_37a2cec8),
    .b(al_bd9d7d67),
    .c(al_f49992c3),
    .o(al_c46301d));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    al_e0ff24b8 (
    .a(al_2c3e73df),
    .b(al_7a486383),
    .c(al_a2deaa78),
    .o(al_f76e538f));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    al_72851dd2 (
    .a(al_6a0e908c),
    .b(al_f76e538f),
    .c(al_6ec8afa5),
    .d(al_a5849610),
    .e(al_e379ebb5),
    .o(al_b279136c));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_ae06f489 (
    .a(al_acd38e8e),
    .b(al_d518b626),
    .o(al_e0005a94));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(C*B))*~(~D*A))"),
    .INIT(32'hff55c040))
    al_734afa27 (
    .a(al_1d3bfd2e),
    .b(al_b279136c),
    .c(al_a8151162),
    .d(al_37a2cec8),
    .e(al_e0005a94),
    .o(al_523a156f));
  AL_MAP_LUT6 #(
    .EQN("(~(F*E*D)*~(A*~(~C*~B)))"),
    .INIT(64'h0057575757575757))
    al_54c42cc2 (
    .a(al_69807e37),
    .b(al_f49992c3),
    .c(al_c73c0ba3),
    .d(al_9b5530fd[0]),
    .e(al_9b5530fd[1]),
    .f(al_9b5530fd[2]),
    .o(al_6e8514b8));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_46dd59e4 (
    .a(al_6e8514b8),
    .b(al_d508bbc9),
    .c(al_6499e5fd),
    .d(al_6893b11d),
    .e(al_f0ecd262),
    .o(al_6a6f79fc));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*A*~(C*B))"),
    .INIT(64'h0000000000002a00))
    al_68c1c690 (
    .a(al_9d63e9cd),
    .b(al_6a0e908c),
    .c(al_5e60a110),
    .d(al_6a6f79fc),
    .e(al_6ec8afa5),
    .f(al_48d2ef94),
    .o(al_7daf5294));
  AL_MAP_LUT6 #(
    .EQN("(~E*B*A*~(C*~(~F*D)))"),
    .INIT(64'h0000080800008808))
    al_c27df997 (
    .a(al_a7b01c14[2]),
    .b(al_7daf5294),
    .c(al_c795a432),
    .d(al_a8151162),
    .e(al_c46301d),
    .f(al_7d2c853e),
    .o(al_cc4ef047));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    al_dfb213c2 (
    .a(al_cc4ef047),
    .b(al_523a156f),
    .c(al_9b5530fd[0]),
    .o(al_c3eb1e82[0]));
  AL_MAP_LUT4 #(
    .EQN("(D@(~(A)*~(B)*~(C)+A*B*C))"),
    .INIT(16'h7e81))
    al_e64dc6d8 (
    .a(al_cc4ef047),
    .b(al_523a156f),
    .c(al_9b5530fd[0]),
    .d(al_9b5530fd[1]),
    .o(al_c3eb1e82[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hdffe8001))
    al_24ebd8f (
    .a(al_cc4ef047),
    .b(al_523a156f),
    .c(al_9b5530fd[0]),
    .d(al_9b5530fd[1]),
    .e(al_9b5530fd[2]),
    .o(al_c3eb1e82[2]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_671640a5 (
    .a(dBusAhb_HREADY_OUT),
    .b(al_aabf3e05),
    .o(dBusAhb_HREADY_IN));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9abdb50a (
    .a(iBusAhb_HRDATA[16]),
    .b(al_b86dd14b[17]),
    .c(al_d518b626),
    .o(al_cf18c1c6[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_691b5df0 (
    .a(iBusAhb_HRDATA[17]),
    .b(al_b86dd14b[18]),
    .c(al_d518b626),
    .o(al_cf18c1c6[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_89b23266 (
    .a(al_b2739b77),
    .b(al_9526c852),
    .c(al_501dbbdf),
    .o(al_a430e4d2));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_420208be (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[5]),
    .o(al_de0f70d9));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_81bdf359 (
    .a(al_85a2bdb0[7]),
    .b(al_85a2bdb0[8]),
    .c(al_85a2bdb0[9]),
    .d(al_85a2bdb0[10]),
    .e(al_85a2bdb0[11]),
    .o(al_1a551855));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hca0fca00))
    al_3c2b959c (
    .a(al_9bcd349b),
    .b(al_e03b3126[16]),
    .c(al_555b0990[0]),
    .d(al_555b0990[1]),
    .e(al_512b1421),
    .o(al_18077581[1]));
  AL_MAP_LUT4 #(
    .EQN("(A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*C*D)"),
    .INIT(16'h8380))
    al_f1a1b6ab (
    .a(al_e03b3126[15]),
    .b(al_555b0990[0]),
    .c(al_555b0990[1]),
    .d(al_1891b3c7),
    .o(al_18077581[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_83c732a5 (
    .a(iBusAhb_HREADY),
    .b(al_a4f21dd7),
    .o(al_acd38e8e));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_344bea2 (
    .a(al_18077581[1]),
    .b(al_2cbb16b4[1]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_201a8a04 (
    .a(al_85a2bdb0[3]),
    .b(al_85a2bdb0[4]),
    .c(al_85a2bdb0[6]),
    .o(al_40a6f08c[29]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_5d980eae (
    .a(al_85a2bdb0[2]),
    .b(al_85a2bdb0[3]),
    .c(al_85a2bdb0[4]),
    .d(al_85a2bdb0[6]),
    .o(al_40a6f08c[30]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_abb0304d (
    .a(al_85a2bdb0[12]),
    .b(al_85a2bdb0[13]),
    .o(al_8bea08a7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f5533000f5533ff))
    al_bc663efc (
    .a(al_e03b3126[7]),
    .b(al_e03b3126[20]),
    .c(al_9bf95cff[0]),
    .d(al_a1e88c0c[0]),
    .e(al_a1e88c0c[1]),
    .f(al_f4b5275b),
    .o(al_f2330f79[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*~A))"),
    .INIT(8'hc9))
    al_19daf261 (
    .a(al_f2330f79[0]),
    .b(al_18077581[0]),
    .c(al_36962d69),
    .o(dBusAhb_HADDR[0]));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*~(C*~(~B*~A)))"),
    .INIT(64'h00001f0000000000))
    al_503ae1a7 (
    .a(dBusAhb_HREADY_OUT),
    .b(al_aabf3e05),
    .c(al_d020f13b),
    .d(al_e3edcf1a),
    .e(al_587b9831),
    .f(al_501dbbdf),
    .o(al_1d840c32));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_6ba9bd62 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .o(al_bb0cd305));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_a0c747ec (
    .a(al_cbdc72d2),
    .b(al_523cde28),
    .o(al_e4d248a4));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0ea0))
    al_92b16b18 (
    .a(dBusAhb_HADDR[0]),
    .b(dBusAhb_HADDR[1]),
    .c(al_bb6625de[1]),
    .d(dBusAhb_HSIZE[1]),
    .o(al_7bc36116));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*~C*~B*~A)"),
    .INIT(64'h0000000001000000))
    al_65a63cb0 (
    .a(al_b469f7cc),
    .b(al_d508bbc9),
    .c(al_6499e5fd),
    .d(al_b567677b),
    .e(al_2a43721c),
    .f(al_6893b11d),
    .o(al_e9d567fe));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_30b1bafb (
    .a(al_e9d567fe),
    .b(al_69807e37),
    .o(al_bec39e4d));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_4878af10 (
    .a(al_e4d248a4),
    .b(al_501dbbdf),
    .c(al_c0a7a5f),
    .o(al_e379ebb5));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h62))
    al_b2f7a712 (
    .a(al_40a6f08c[30]),
    .b(al_40a6f08c[29]),
    .c(al_85a2bdb0[31]),
    .o(al_da9c21fb));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    al_576820d0 (
    .a(al_c73c0ba3),
    .b(al_5c72a609[1]),
    .c(al_5c72a609[2]),
    .o(al_f6cd735f));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_d312dd6f (
    .a(al_8bf5da64),
    .b(al_523cde28),
    .o(al_b211b12d));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_75c32e1d (
    .a(al_bec39e4d),
    .b(al_5e275e81),
    .o(al_c91705db));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_9315568c (
    .a(al_212ac3ba[0]),
    .b(al_212ac3ba[1]),
    .c(al_c0a7a5f),
    .o(al_ea2eaeb1));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_2e939c4b (
    .a(al_c91705db),
    .b(al_ea2eaeb1),
    .o(al_9d63e9cd));
  AL_MAP_LUT6 #(
    .EQN("(~E*~(~F*D*~C*B*A))"),
    .INIT(64'h0000ffff0000f7ff))
    al_1e002977 (
    .a(dBusAhb_HREADY_OUT),
    .b(dBusAhb_HRESP),
    .c(al_aabf3e05),
    .d(al_d020f13b),
    .e(al_673a4598),
    .f(al_587b9831),
    .o(al_68b106c6));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_962c8674 (
    .a(al_68b106c6),
    .b(al_e3edcf1a),
    .c(al_501dbbdf),
    .o(al_6ec8afa5));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_7867816c (
    .a(al_202f2c67[0]),
    .b(al_202f2c67[1]),
    .c(al_202f2c67[2]),
    .o(al_7a486383));
  AL_MAP_LUT6 #(
    .EQN("(D*A*~(~(~C*B)*~(E)*~(F)+~(~C*B)*E*~(F)+~(~(~C*B))*E*F+~(~C*B)*E*F))"),
    .INIT(64'h0000aa0008000800))
    al_54115ddd (
    .a(al_7a486383),
    .b(al_acd38e8e),
    .c(iBusAhb_HRESP),
    .d(al_f49992c3),
    .e(al_b86dd14b[0]),
    .f(al_d518b626),
    .o(al_bd9d7d67));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_aa64a756 (
    .a(al_85a2bdb0[20]),
    .b(al_85a2bdb0[21]),
    .c(al_85a2bdb0[23]),
    .d(al_a0e6869c[7]),
    .e(al_a0e6869c[8]),
    .f(al_a0e6869c[10]),
    .o(al_2f23ede9));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_fecb3245 (
    .a(al_2f23ede9),
    .b(al_85a2bdb0[22]),
    .c(al_85a2bdb0[24]),
    .d(al_a0e6869c[9]),
    .e(al_a0e6869c[11]),
    .o(al_df2df2f9));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_44ead8a8 (
    .a(al_85a2bdb0[20]),
    .b(al_85a2bdb0[21]),
    .c(al_85a2bdb0[22]),
    .d(al_e03b3126[7]),
    .e(al_e03b3126[8]),
    .f(al_e03b3126[9]),
    .o(al_689ac380));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_d1ea4953 (
    .a(al_689ac380),
    .b(al_85a2bdb0[23]),
    .c(al_85a2bdb0[24]),
    .d(al_e03b3126[10]),
    .e(al_e03b3126[11]),
    .o(al_358f5bea));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_a0aecb68 (
    .a(al_85a2bdb0[15]),
    .b(al_85a2bdb0[16]),
    .c(al_85a2bdb0[18]),
    .d(al_a0e6869c[7]),
    .e(al_a0e6869c[8]),
    .f(al_a0e6869c[10]),
    .o(al_17050ddb));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_f208f711 (
    .a(al_17050ddb),
    .b(al_85a2bdb0[17]),
    .c(al_85a2bdb0[19]),
    .d(al_a0e6869c[9]),
    .e(al_a0e6869c[11]),
    .o(al_a2426a1));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_7994955d (
    .a(al_85a2bdb0[15]),
    .b(al_85a2bdb0[16]),
    .c(al_85a2bdb0[17]),
    .d(al_e03b3126[7]),
    .e(al_e03b3126[8]),
    .f(al_e03b3126[9]),
    .o(al_6faa66d6));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_34c4c48c (
    .a(al_3ca44efd[0]),
    .o({al_e9183b70,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_799b81f8 (
    .a(al_df7b4407),
    .b(al_18077581[0]),
    .c(al_e9183b70),
    .o({al_7709e0b8,open_n23}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_95a9b52b (
    .a(al_18077581[1]),
    .b(al_3ca44efd[1]),
    .c(al_7709e0b8),
    .o({al_5907d462,al_2cbb16b4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_852c4c0c (
    .a(al_18077581[2]),
    .b(al_3ca44efd[2]),
    .c(al_5907d462),
    .o({al_e83c9381,al_2cbb16b4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4e157650 (
    .a(al_18077581[3]),
    .b(al_3ca44efd[3]),
    .c(al_e83c9381),
    .o({al_b4c2dbf,al_2cbb16b4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1f3a8851 (
    .a(al_18077581[4]),
    .b(al_3ca44efd[4]),
    .c(al_b4c2dbf),
    .o({al_cd728703,al_2cbb16b4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_524b4e57 (
    .a(al_18077581[5]),
    .b(al_3ca44efd[5]),
    .c(al_cd728703),
    .o({al_6dc2ee9d,al_2cbb16b4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3dab8fb8 (
    .a(al_18077581[6]),
    .b(al_3ca44efd[6]),
    .c(al_6dc2ee9d),
    .o({al_36d94dee,al_2cbb16b4[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_33929a09 (
    .a(al_18077581[7]),
    .b(al_3ca44efd[7]),
    .c(al_36d94dee),
    .o({al_e493cfe2,al_2cbb16b4[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d3c59aaf (
    .a(al_18077581[8]),
    .b(al_3ca44efd[8]),
    .c(al_e493cfe2),
    .o({al_a122473,al_2cbb16b4[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_708c43c4 (
    .a(al_18077581[9]),
    .b(al_3ca44efd[9]),
    .c(al_a122473),
    .o({al_571b50e9,al_2cbb16b4[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4978b26a (
    .a(al_18077581[10]),
    .b(al_3ca44efd[10]),
    .c(al_571b50e9),
    .o({al_91e1bb2e,al_2cbb16b4[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_485e77ec (
    .a(al_18077581[11]),
    .b(al_3ca44efd[11]),
    .c(al_91e1bb2e),
    .o({al_89941f61,al_2cbb16b4[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3b06e2f7 (
    .a(al_18077581[12]),
    .b(al_3ca44efd[12]),
    .c(al_89941f61),
    .o({al_57355198,al_2cbb16b4[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a6cb7175 (
    .a(al_18077581[13]),
    .b(al_3ca44efd[13]),
    .c(al_57355198),
    .o({al_c768664c,al_2cbb16b4[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b5dcd95e (
    .a(al_18077581[14]),
    .b(al_3ca44efd[14]),
    .c(al_c768664c),
    .o({al_7e44038b,al_2cbb16b4[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ddaf73df (
    .a(al_18077581[15]),
    .b(al_3ca44efd[15]),
    .c(al_7e44038b),
    .o({al_c6e3e50,al_2cbb16b4[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b088bd8a (
    .a(al_18077581[16]),
    .b(al_3ca44efd[16]),
    .c(al_c6e3e50),
    .o({al_58a3b7ac,al_2cbb16b4[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9b7e6b9c (
    .a(al_18077581[17]),
    .b(al_3ca44efd[17]),
    .c(al_58a3b7ac),
    .o({al_fe608411,al_2cbb16b4[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1a1d1fb3 (
    .a(al_18077581[18]),
    .b(al_3ca44efd[18]),
    .c(al_fe608411),
    .o({al_a8c327eb,al_2cbb16b4[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_73082578 (
    .a(al_18077581[19]),
    .b(al_3ca44efd[19]),
    .c(al_a8c327eb),
    .o({al_c02355f,al_2cbb16b4[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3759d498 (
    .a(al_18077581[20]),
    .b(al_3ca44efd[20]),
    .c(al_c02355f),
    .o({al_50f055e6,al_2cbb16b4[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f67b37dc (
    .a(al_18077581[21]),
    .b(al_3ca44efd[21]),
    .c(al_50f055e6),
    .o({al_7971debc,al_2cbb16b4[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5097520c (
    .a(al_18077581[22]),
    .b(al_3ca44efd[22]),
    .c(al_7971debc),
    .o({al_8628bcb0,al_2cbb16b4[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cf6a99db (
    .a(al_18077581[23]),
    .b(al_3ca44efd[23]),
    .c(al_8628bcb0),
    .o({al_5d524bff,al_2cbb16b4[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_68bfea03 (
    .a(al_18077581[24]),
    .b(al_3ca44efd[24]),
    .c(al_5d524bff),
    .o({al_ed4da032,al_2cbb16b4[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_924f197f (
    .a(al_18077581[25]),
    .b(al_3ca44efd[25]),
    .c(al_ed4da032),
    .o({al_931aa04b,al_2cbb16b4[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_620ced48 (
    .a(al_18077581[26]),
    .b(al_3ca44efd[26]),
    .c(al_931aa04b),
    .o({al_571c1ade,al_2cbb16b4[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9796fb79 (
    .a(al_18077581[27]),
    .b(al_3ca44efd[27]),
    .c(al_571c1ade),
    .o({al_7d44614a,al_2cbb16b4[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c91059a2 (
    .a(al_18077581[28]),
    .b(al_3ca44efd[28]),
    .c(al_7d44614a),
    .o({al_fc020630,al_2cbb16b4[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_db5299f4 (
    .a(al_18077581[29]),
    .b(al_3ca44efd[29]),
    .c(al_fc020630),
    .o({al_381491bf,al_2cbb16b4[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ff829624 (
    .a(al_18077581[30]),
    .b(al_3ca44efd[30]),
    .c(al_381491bf),
    .o({al_862095a3,al_2cbb16b4[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f6373967 (
    .a(al_18077581[31]),
    .b(al_3ca44efd[31]),
    .c(al_862095a3),
    .o({open_n24,al_2cbb16b4[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_aea212eb (
    .a(1'b0),
    .o({al_d81efc87,open_n27}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_63be8699 (
    .a(al_f3b8f942[0]),
    .b(al_a167c8cf),
    .c(al_d81efc87),
    .o({al_afa2ef7a,open_n28}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a7ad2865 (
    .a(al_f3b8f942[1]),
    .b(1'b0),
    .c(al_afa2ef7a),
    .o({al_5a473143,al_32172a12[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1833fd92 (
    .a(al_f3b8f942[2]),
    .b(1'b0),
    .c(al_5a473143),
    .o({al_9a380597,al_32172a12[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a3a39408 (
    .a(al_f3b8f942[3]),
    .b(1'b0),
    .c(al_9a380597),
    .o({al_2fd5db25,al_32172a12[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9bed92dc (
    .a(al_f3b8f942[4]),
    .b(1'b0),
    .c(al_2fd5db25),
    .o({al_83abb1fc,al_32172a12[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4d6b5b0a (
    .a(al_f3b8f942[5]),
    .b(1'b0),
    .c(al_83abb1fc),
    .o({al_bb6e1564,al_32172a12[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d32e784a (
    .a(al_f3b8f942[6]),
    .b(1'b0),
    .c(al_bb6e1564),
    .o({al_76d86d60,al_32172a12[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_92f7d7f0 (
    .a(al_f3b8f942[7]),
    .b(1'b0),
    .c(al_76d86d60),
    .o({al_abafb840,al_32172a12[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_424ee8c9 (
    .a(al_f3b8f942[8]),
    .b(1'b0),
    .c(al_abafb840),
    .o({al_665b60c1,al_32172a12[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8f962df (
    .a(al_f3b8f942[9]),
    .b(1'b0),
    .c(al_665b60c1),
    .o({al_9367b2dc,al_32172a12[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_48397d16 (
    .a(al_f3b8f942[10]),
    .b(1'b0),
    .c(al_9367b2dc),
    .o({al_e6c5dfa,al_32172a12[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b2cb5b29 (
    .a(al_f3b8f942[11]),
    .b(1'b0),
    .c(al_e6c5dfa),
    .o({al_5188e109,al_32172a12[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8f3fdd08 (
    .a(al_f3b8f942[12]),
    .b(1'b0),
    .c(al_5188e109),
    .o({al_75b52645,al_32172a12[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b7743a27 (
    .a(al_f3b8f942[13]),
    .b(1'b0),
    .c(al_75b52645),
    .o({al_20769005,al_32172a12[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b6cba910 (
    .a(al_f3b8f942[14]),
    .b(1'b0),
    .c(al_20769005),
    .o({al_4d3a4f57,al_32172a12[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ef69e78d (
    .a(al_f3b8f942[15]),
    .b(1'b0),
    .c(al_4d3a4f57),
    .o({al_ead254a9,al_32172a12[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1d2b030 (
    .a(al_f3b8f942[16]),
    .b(1'b0),
    .c(al_ead254a9),
    .o({al_bdce010d,al_32172a12[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d4007e82 (
    .a(al_f3b8f942[17]),
    .b(1'b0),
    .c(al_bdce010d),
    .o({al_8cc085cf,al_32172a12[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_703012d8 (
    .a(al_f3b8f942[18]),
    .b(1'b0),
    .c(al_8cc085cf),
    .o({al_83e5bc67,al_32172a12[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e5f70ffc (
    .a(al_f3b8f942[19]),
    .b(1'b0),
    .c(al_83e5bc67),
    .o({al_cc21f874,al_32172a12[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d7531e6c (
    .a(al_f3b8f942[20]),
    .b(1'b0),
    .c(al_cc21f874),
    .o({al_304a2593,al_32172a12[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c900c823 (
    .a(al_f3b8f942[21]),
    .b(1'b0),
    .c(al_304a2593),
    .o({al_de514d5,al_32172a12[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_81d2247f (
    .a(al_f3b8f942[22]),
    .b(1'b0),
    .c(al_de514d5),
    .o({al_3178c29a,al_32172a12[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_95237b75 (
    .a(al_f3b8f942[23]),
    .b(1'b0),
    .c(al_3178c29a),
    .o({al_bf8b5005,al_32172a12[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_612e5f34 (
    .a(al_f3b8f942[24]),
    .b(1'b0),
    .c(al_bf8b5005),
    .o({al_322e0ef8,al_32172a12[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1c0a6cd5 (
    .a(al_f3b8f942[25]),
    .b(1'b0),
    .c(al_322e0ef8),
    .o({al_9cc77063,al_32172a12[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_46c4c171 (
    .a(al_f3b8f942[26]),
    .b(1'b0),
    .c(al_9cc77063),
    .o({al_5c37ca50,al_32172a12[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_48dc238 (
    .a(al_f3b8f942[27]),
    .b(1'b0),
    .c(al_5c37ca50),
    .o({al_7e8c6cca,al_32172a12[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6c689a0b (
    .a(al_f3b8f942[28]),
    .b(1'b0),
    .c(al_7e8c6cca),
    .o({al_1b896d0b,al_32172a12[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b3b0e45 (
    .a(al_f3b8f942[29]),
    .b(1'b0),
    .c(al_1b896d0b),
    .o({al_a8c77bd0,al_32172a12[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_daf73106 (
    .a(al_f3b8f942[30]),
    .b(1'b0),
    .c(al_a8c77bd0),
    .o({al_3d1aa152,al_32172a12[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c5392032 (
    .a(al_f3b8f942[31]),
    .b(1'b0),
    .c(al_3d1aa152),
    .o({open_n29,al_32172a12[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_3abc2cff (
    .a(1'b0),
    .o({al_3c0b578d,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b233958a (
    .a(al_d57349d9[0]),
    .b(al_35295e0a[0]),
    .c(al_3c0b578d),
    .o({al_8c1979b0,open_n33}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3f25f89c (
    .a(al_d57349d9[1]),
    .b(al_35295e0a[1]),
    .c(al_8c1979b0),
    .o({al_6a1d2e79,al_6f2fa5dc[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4725daf5 (
    .a(al_d57349d9[2]),
    .b(al_35295e0a[2]),
    .c(al_6a1d2e79),
    .o({al_1520e815,al_6f2fa5dc[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dc083b74 (
    .a(al_d57349d9[3]),
    .b(al_35295e0a[3]),
    .c(al_1520e815),
    .o({al_7bc70fec,al_6f2fa5dc[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b5f7a822 (
    .a(al_d57349d9[4]),
    .b(al_35295e0a[4]),
    .c(al_7bc70fec),
    .o({al_5b63e1bd,al_6f2fa5dc[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7e989d87 (
    .a(al_d57349d9[5]),
    .b(al_35295e0a[5]),
    .c(al_5b63e1bd),
    .o({al_c30b4452,al_6f2fa5dc[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_40e170dc (
    .a(al_d57349d9[6]),
    .b(al_35295e0a[6]),
    .c(al_c30b4452),
    .o({al_1da1b47c,al_6f2fa5dc[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b2f4a043 (
    .a(al_d57349d9[7]),
    .b(al_35295e0a[7]),
    .c(al_1da1b47c),
    .o({al_f380f225,al_6f2fa5dc[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_45fef5ec (
    .a(al_d57349d9[8]),
    .b(al_35295e0a[8]),
    .c(al_f380f225),
    .o({al_c45763da,al_6f2fa5dc[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ed5ee606 (
    .a(al_d57349d9[9]),
    .b(al_35295e0a[9]),
    .c(al_c45763da),
    .o({al_91dd025b,al_6f2fa5dc[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_447df3da (
    .a(al_d57349d9[10]),
    .b(al_35295e0a[10]),
    .c(al_91dd025b),
    .o({al_1e473c0d,al_6f2fa5dc[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_841d4a30 (
    .a(al_d57349d9[11]),
    .b(al_35295e0a[11]),
    .c(al_1e473c0d),
    .o({al_429b8bb,al_6f2fa5dc[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f9d223d7 (
    .a(al_d57349d9[12]),
    .b(al_35295e0a[12]),
    .c(al_429b8bb),
    .o({al_a0d06894,al_6f2fa5dc[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ce0b130d (
    .a(al_d57349d9[13]),
    .b(al_35295e0a[13]),
    .c(al_a0d06894),
    .o({al_ab3758ac,al_6f2fa5dc[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c244238b (
    .a(al_d57349d9[14]),
    .b(al_35295e0a[14]),
    .c(al_ab3758ac),
    .o({al_399d7ca4,al_6f2fa5dc[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e715d7c0 (
    .a(al_d57349d9[15]),
    .b(al_35295e0a[15]),
    .c(al_399d7ca4),
    .o({al_e87887db,al_6f2fa5dc[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_59021e55 (
    .a(al_d57349d9[16]),
    .b(al_35295e0a[16]),
    .c(al_e87887db),
    .o({al_252ad8ef,al_6f2fa5dc[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_906b7510 (
    .a(al_d57349d9[17]),
    .b(al_35295e0a[17]),
    .c(al_252ad8ef),
    .o({al_ed00e897,al_6f2fa5dc[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a8c57bc4 (
    .a(al_d57349d9[18]),
    .b(al_35295e0a[18]),
    .c(al_ed00e897),
    .o({al_5ab03ac,al_6f2fa5dc[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bb16147a (
    .a(al_d57349d9[19]),
    .b(al_35295e0a[19]),
    .c(al_5ab03ac),
    .o({al_6afd474a,al_6f2fa5dc[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_40c5d44 (
    .a(al_d57349d9[20]),
    .b(al_35295e0a[20]),
    .c(al_6afd474a),
    .o({al_ae709366,al_6f2fa5dc[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_68db6e13 (
    .a(al_d57349d9[21]),
    .b(al_35295e0a[20]),
    .c(al_ae709366),
    .o({al_1a6b06a2,al_6f2fa5dc[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c92360e9 (
    .a(al_d57349d9[22]),
    .b(al_35295e0a[20]),
    .c(al_1a6b06a2),
    .o({al_630fb1c3,al_6f2fa5dc[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c50aa0a2 (
    .a(al_d57349d9[23]),
    .b(al_35295e0a[20]),
    .c(al_630fb1c3),
    .o({al_ac5e9239,al_6f2fa5dc[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e1cb90a8 (
    .a(al_d57349d9[24]),
    .b(al_35295e0a[20]),
    .c(al_ac5e9239),
    .o({al_f58e845f,al_6f2fa5dc[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_69685ad5 (
    .a(al_d57349d9[25]),
    .b(al_35295e0a[20]),
    .c(al_f58e845f),
    .o({al_388498bb,al_6f2fa5dc[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_42e63541 (
    .a(al_d57349d9[26]),
    .b(al_35295e0a[20]),
    .c(al_388498bb),
    .o({al_9ef79df4,al_6f2fa5dc[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_35b7a39a (
    .a(al_d57349d9[27]),
    .b(al_35295e0a[20]),
    .c(al_9ef79df4),
    .o({al_818b914,al_6f2fa5dc[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1421b73e (
    .a(al_d57349d9[28]),
    .b(al_35295e0a[20]),
    .c(al_818b914),
    .o({al_b113fb3b,al_6f2fa5dc[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b90ec81a (
    .a(al_d57349d9[29]),
    .b(al_35295e0a[20]),
    .c(al_b113fb3b),
    .o({al_614db1c3,al_6f2fa5dc[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_398dc396 (
    .a(al_d57349d9[30]),
    .b(al_35295e0a[20]),
    .c(al_614db1c3),
    .o({al_8dd6f665,al_6f2fa5dc[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d218e0e7 (
    .a(al_d57349d9[31]),
    .b(al_35295e0a[20]),
    .c(al_8dd6f665),
    .o({open_n34,al_6f2fa5dc[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_67457eb7 (
    .a(1'b0),
    .o({al_2340ada,open_n37}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a7aa3552 (
    .a(al_439698e9[0]),
    .b(al_698ba8c2),
    .c(al_2340ada),
    .o({al_6233890d,open_n38}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_37626348 (
    .a(al_439698e9[1]),
    .b(1'b0),
    .c(al_6233890d),
    .o({al_d0d487f0,al_afda7fe3[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b8883486 (
    .a(al_439698e9[2]),
    .b(1'b0),
    .c(al_d0d487f0),
    .o({al_f5ef5e84,al_afda7fe3[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_abf2597a (
    .a(al_439698e9[3]),
    .b(1'b0),
    .c(al_f5ef5e84),
    .o({al_dea86dcd,al_afda7fe3[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e2506647 (
    .a(al_439698e9[4]),
    .b(1'b0),
    .c(al_dea86dcd),
    .o({al_429d51be,al_afda7fe3[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_865ca757 (
    .a(al_439698e9[5]),
    .b(1'b0),
    .c(al_429d51be),
    .o({al_c5f16127,al_afda7fe3[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_40f98bfa (
    .a(al_439698e9[6]),
    .b(1'b0),
    .c(al_c5f16127),
    .o({al_9b8294d5,al_afda7fe3[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_adcc35ea (
    .a(al_439698e9[7]),
    .b(1'b0),
    .c(al_9b8294d5),
    .o({al_382bcd96,al_afda7fe3[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_54f748f7 (
    .a(al_439698e9[8]),
    .b(1'b0),
    .c(al_382bcd96),
    .o({al_59258acc,al_afda7fe3[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d517902c (
    .a(al_439698e9[9]),
    .b(1'b0),
    .c(al_59258acc),
    .o({al_5a3cd9,al_afda7fe3[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_48ba439d (
    .a(al_439698e9[10]),
    .b(1'b0),
    .c(al_5a3cd9),
    .o({al_e3fa7139,al_afda7fe3[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1805ef5b (
    .a(al_439698e9[11]),
    .b(1'b0),
    .c(al_e3fa7139),
    .o({al_a4b5d1d0,al_afda7fe3[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_30dafe3 (
    .a(al_439698e9[12]),
    .b(1'b0),
    .c(al_a4b5d1d0),
    .o({al_774d209c,al_afda7fe3[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e31c315b (
    .a(al_439698e9[13]),
    .b(1'b0),
    .c(al_774d209c),
    .o({al_eecd0df4,al_afda7fe3[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_810efd57 (
    .a(al_439698e9[14]),
    .b(1'b0),
    .c(al_eecd0df4),
    .o({al_491245fc,al_afda7fe3[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cc600473 (
    .a(al_439698e9[15]),
    .b(1'b0),
    .c(al_491245fc),
    .o({al_151b9283,al_afda7fe3[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a489f7c6 (
    .a(al_439698e9[16]),
    .b(1'b0),
    .c(al_151b9283),
    .o({al_aac49860,al_afda7fe3[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_81f79c52 (
    .a(al_439698e9[17]),
    .b(1'b0),
    .c(al_aac49860),
    .o({al_826899ea,al_afda7fe3[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_606a06b2 (
    .a(al_439698e9[18]),
    .b(1'b0),
    .c(al_826899ea),
    .o({al_3401493,al_afda7fe3[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_303411a7 (
    .a(al_439698e9[19]),
    .b(1'b0),
    .c(al_3401493),
    .o({al_e381eae8,al_afda7fe3[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_71f94044 (
    .a(al_439698e9[20]),
    .b(1'b0),
    .c(al_e381eae8),
    .o({al_29590532,al_afda7fe3[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d680521c (
    .a(al_439698e9[21]),
    .b(1'b0),
    .c(al_29590532),
    .o({al_a5dcf577,al_afda7fe3[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_90ebec12 (
    .a(al_439698e9[22]),
    .b(1'b0),
    .c(al_a5dcf577),
    .o({al_f20e1999,al_afda7fe3[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b73afe58 (
    .a(al_439698e9[23]),
    .b(1'b0),
    .c(al_f20e1999),
    .o({al_9f91dd62,al_afda7fe3[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3f66d5da (
    .a(al_439698e9[24]),
    .b(1'b0),
    .c(al_9f91dd62),
    .o({al_4945d0da,al_afda7fe3[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_417cb907 (
    .a(al_439698e9[25]),
    .b(1'b0),
    .c(al_4945d0da),
    .o({al_7cba307c,al_afda7fe3[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2238c9ca (
    .a(al_439698e9[26]),
    .b(1'b0),
    .c(al_7cba307c),
    .o({al_50fdf48e,al_afda7fe3[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2d500183 (
    .a(al_439698e9[27]),
    .b(1'b0),
    .c(al_50fdf48e),
    .o({al_bc2094a,al_afda7fe3[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_43281ae (
    .a(al_439698e9[28]),
    .b(1'b0),
    .c(al_bc2094a),
    .o({al_be7d7ec3,al_afda7fe3[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6a36165e (
    .a(al_439698e9[29]),
    .b(1'b0),
    .c(al_be7d7ec3),
    .o({al_7c4abb1c,al_afda7fe3[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1d5365bd (
    .a(al_439698e9[30]),
    .b(1'b0),
    .c(al_7c4abb1c),
    .o({al_35216c23,al_afda7fe3[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_629e92bf (
    .a(al_439698e9[31]),
    .b(1'b0),
    .c(al_35216c23),
    .o({open_n39,al_afda7fe3[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_51a12919 (
    .a(1'b0),
    .o({al_34eb7e40,open_n42}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_562e45cf (
    .a(al_4e7a070d[0]),
    .b(al_ba08f61a),
    .c(al_34eb7e40),
    .o({al_8bbc936e,open_n43}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_155b727c (
    .a(al_4e7a070d[1]),
    .b(1'b0),
    .c(al_8bbc936e),
    .o({al_33f7e9f,al_f337bb3c[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4e486993 (
    .a(al_4e7a070d[2]),
    .b(1'b0),
    .c(al_33f7e9f),
    .o({al_82cf60b4,al_f337bb3c[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_694186b8 (
    .a(al_4e7a070d[3]),
    .b(1'b0),
    .c(al_82cf60b4),
    .o({al_87a252af,al_f337bb3c[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_75152959 (
    .a(al_4e7a070d[4]),
    .b(1'b0),
    .c(al_87a252af),
    .o({al_e2de4855,al_f337bb3c[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2cfb7b5c (
    .a(al_4e7a070d[5]),
    .b(1'b0),
    .c(al_e2de4855),
    .o({al_6e34d4cd,al_f337bb3c[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cca81331 (
    .a(al_4e7a070d[6]),
    .b(1'b0),
    .c(al_6e34d4cd),
    .o({al_1af3cc59,al_f337bb3c[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_40662957 (
    .a(al_4e7a070d[7]),
    .b(1'b0),
    .c(al_1af3cc59),
    .o({al_2161900e,al_f337bb3c[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6c5e729 (
    .a(al_4e7a070d[8]),
    .b(1'b0),
    .c(al_2161900e),
    .o({al_eba13280,al_f337bb3c[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c0898dca (
    .a(al_4e7a070d[9]),
    .b(1'b0),
    .c(al_eba13280),
    .o({al_837ccd29,al_f337bb3c[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_301b2a24 (
    .a(al_4e7a070d[10]),
    .b(1'b0),
    .c(al_837ccd29),
    .o({al_9711882c,al_f337bb3c[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a55d4bf2 (
    .a(al_4e7a070d[11]),
    .b(1'b0),
    .c(al_9711882c),
    .o({al_2d65cded,al_f337bb3c[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6056132f (
    .a(al_4e7a070d[12]),
    .b(1'b0),
    .c(al_2d65cded),
    .o({al_de77c599,al_f337bb3c[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_55cf1325 (
    .a(al_4e7a070d[13]),
    .b(1'b0),
    .c(al_de77c599),
    .o({al_e2f41361,al_f337bb3c[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5af9da00 (
    .a(al_4e7a070d[14]),
    .b(1'b0),
    .c(al_e2f41361),
    .o({al_af2b71d8,al_f337bb3c[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7de456e3 (
    .a(al_4e7a070d[15]),
    .b(1'b0),
    .c(al_af2b71d8),
    .o({al_96191e5,al_f337bb3c[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7376fe0e (
    .a(al_4e7a070d[16]),
    .b(1'b0),
    .c(al_96191e5),
    .o({al_b81cc851,al_f337bb3c[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2f14a033 (
    .a(al_4e7a070d[17]),
    .b(1'b0),
    .c(al_b81cc851),
    .o({al_1af8f97e,al_f337bb3c[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fc0ec398 (
    .a(al_4e7a070d[18]),
    .b(1'b0),
    .c(al_1af8f97e),
    .o({al_4db67ec5,al_f337bb3c[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b8f73752 (
    .a(al_4e7a070d[19]),
    .b(1'b0),
    .c(al_4db67ec5),
    .o({al_24887a1a,al_f337bb3c[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_559a5ec3 (
    .a(al_4e7a070d[20]),
    .b(1'b0),
    .c(al_24887a1a),
    .o({al_9a21e871,al_f337bb3c[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_de83172b (
    .a(al_4e7a070d[21]),
    .b(1'b0),
    .c(al_9a21e871),
    .o({al_35d69006,al_f337bb3c[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6057c5c8 (
    .a(al_4e7a070d[22]),
    .b(1'b0),
    .c(al_35d69006),
    .o({al_d3f03020,al_f337bb3c[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_91866ae (
    .a(al_4e7a070d[23]),
    .b(1'b0),
    .c(al_d3f03020),
    .o({al_2d292595,al_f337bb3c[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2c3730b8 (
    .a(al_4e7a070d[24]),
    .b(1'b0),
    .c(al_2d292595),
    .o({al_5325cd47,al_f337bb3c[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bb0eb211 (
    .a(al_4e7a070d[25]),
    .b(1'b0),
    .c(al_5325cd47),
    .o({al_bf79dcf1,al_f337bb3c[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f5237083 (
    .a(al_4e7a070d[26]),
    .b(1'b0),
    .c(al_bf79dcf1),
    .o({al_58ec462a,al_f337bb3c[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9de53236 (
    .a(al_4e7a070d[27]),
    .b(1'b0),
    .c(al_58ec462a),
    .o({al_42d8598b,al_f337bb3c[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d3a3bf10 (
    .a(al_4e7a070d[28]),
    .b(1'b0),
    .c(al_42d8598b),
    .o({al_9bb4d4a4,al_f337bb3c[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4b81c98e (
    .a(al_4e7a070d[29]),
    .b(1'b0),
    .c(al_9bb4d4a4),
    .o({al_82229532,al_f337bb3c[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1f4a7350 (
    .a(al_4e7a070d[30]),
    .b(1'b0),
    .c(al_82229532),
    .o({al_ec42a4de,al_f337bb3c[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_282752b2 (
    .a(al_4e7a070d[31]),
    .b(1'b0),
    .c(al_ec42a4de),
    .o({open_n44,al_f337bb3c[31]}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_7e95ea91 (
    .a(dBusAhb_HRDATA[0]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[0]),
    .o(al_8c4e5d9c[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_5a817fca (
    .a(dBusAhb_HRDATA[10]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[10]),
    .o(al_8c4e5d9c[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_efac656 (
    .a(dBusAhb_HRDATA[11]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[11]),
    .o(al_8c4e5d9c[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_3d722544 (
    .a(dBusAhb_HRDATA[12]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[12]),
    .o(al_8c4e5d9c[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_841cca07 (
    .a(dBusAhb_HRDATA[13]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[13]),
    .o(al_8c4e5d9c[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_bad960b5 (
    .a(dBusAhb_HRDATA[14]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[14]),
    .o(al_8c4e5d9c[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_851d3441 (
    .a(dBusAhb_HRDATA[15]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[15]),
    .o(al_8c4e5d9c[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_432142a9 (
    .a(dBusAhb_HRDATA[16]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[16]),
    .o(al_8c4e5d9c[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_b6b06e30 (
    .a(dBusAhb_HRDATA[17]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[17]),
    .o(al_8c4e5d9c[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_5be8932c (
    .a(dBusAhb_HRDATA[18]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[18]),
    .o(al_8c4e5d9c[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_84e784c7 (
    .a(dBusAhb_HRDATA[19]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[19]),
    .o(al_8c4e5d9c[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_98640e24 (
    .a(dBusAhb_HRDATA[1]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[1]),
    .o(al_8c4e5d9c[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_6d3b3107 (
    .a(dBusAhb_HRDATA[20]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[20]),
    .o(al_8c4e5d9c[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_c58debd7 (
    .a(dBusAhb_HRDATA[21]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[21]),
    .o(al_8c4e5d9c[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_83c3c0b7 (
    .a(dBusAhb_HRDATA[22]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[22]),
    .o(al_8c4e5d9c[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_57cfa912 (
    .a(dBusAhb_HRDATA[23]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[23]),
    .o(al_8c4e5d9c[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_cb2a101e (
    .a(dBusAhb_HRDATA[24]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[24]),
    .o(al_8c4e5d9c[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_7229c1a1 (
    .a(dBusAhb_HRDATA[25]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[25]),
    .o(al_8c4e5d9c[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_29275b5e (
    .a(dBusAhb_HRDATA[26]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[26]),
    .o(al_8c4e5d9c[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_5d2c2c6b (
    .a(dBusAhb_HRDATA[27]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[27]),
    .o(al_8c4e5d9c[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_ca15ad4b (
    .a(dBusAhb_HRDATA[28]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[28]),
    .o(al_8c4e5d9c[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_9aa5aedd (
    .a(dBusAhb_HRDATA[29]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[29]),
    .o(al_8c4e5d9c[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_128c8f93 (
    .a(dBusAhb_HRDATA[2]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[2]),
    .o(al_8c4e5d9c[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_6e3953f7 (
    .a(dBusAhb_HRDATA[30]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[30]),
    .o(al_8c4e5d9c[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_1b615141 (
    .a(dBusAhb_HRDATA[3]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[3]),
    .o(al_8c4e5d9c[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_7c6d0b62 (
    .a(dBusAhb_HRDATA[4]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[4]),
    .o(al_8c4e5d9c[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_a2ca9c6d (
    .a(dBusAhb_HRDATA[5]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[5]),
    .o(al_8c4e5d9c[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_210d0051 (
    .a(dBusAhb_HRDATA[6]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[6]),
    .o(al_8c4e5d9c[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_27dcf9fd (
    .a(dBusAhb_HRDATA[7]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[7]),
    .o(al_8c4e5d9c[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_86ca42c7 (
    .a(dBusAhb_HRDATA[8]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[8]),
    .o(al_8c4e5d9c[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_427f5dfa (
    .a(dBusAhb_HRDATA[9]),
    .b(al_aabf3e05),
    .c(al_7c5dfaf6[9]),
    .o(al_8c4e5d9c[9]));
  AL_DFF_X al_6971797a (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_681bbb63),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18c565c8));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_452f4956 (
    .a(al_8a4a038[1]),
    .b(al_8a4a038[2]),
    .c(al_8a4a038[3]),
    .d(al_8a4a038[4]),
    .e(al_8a4a038[5]),
    .f(al_8a4a038[6]),
    .o(al_510fa565));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_af5ecba6 (
    .a(al_510fa565),
    .b(al_a7af1013),
    .c(al_8a4a038[0]),
    .d(al_8a4a038[7]),
    .o(al_4cb17b0d));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_26c940f3 (
    .a(al_4cb17b0d),
    .b(al_cb807890),
    .o(al_681bbb63));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_24363fc6 (
    .a(al_1a551855),
    .b(al_85a2bdb0[12]),
    .c(al_85a2bdb0[13]),
    .o(al_566f1754));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~E*~D*~C*~B*A)"),
    .INIT(64'hfffffffffffffffd))
    al_39b48341 (
    .a(al_85a2bdb0[13]),
    .b(al_85a2bdb0[15]),
    .c(al_85a2bdb0[16]),
    .d(al_85a2bdb0[17]),
    .e(al_85a2bdb0[18]),
    .f(al_85a2bdb0[19]),
    .o(al_2434efda));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    al_60f013bb (
    .a(al_8bea08a7),
    .b(al_6893b11d),
    .c(al_85a2bdb0[4]),
    .d(al_85a2bdb0[6]),
    .e(al_85a2bdb0[20]),
    .o(al_5978317));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_bca0e884 (
    .a(al_5978317),
    .b(al_afb86315),
    .c(al_67635cb3),
    .d(al_85a2bdb0[28]),
    .o(al_c4aa9af));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_4722c887 (
    .a(al_fb22b66),
    .b(al_a7b01c14[2]),
    .c(al_85a2bdb0[15]),
    .o(al_704d20e3[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B*~A))"),
    .INIT(8'h4f))
    al_58faa77e (
    .a(al_9ae3000c),
    .b(al_dec34edc),
    .c(al_5c28a20d),
    .o(al_704d20e3[16]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    .INIT(16'hfbc8))
    al_98b0bcfe (
    .a(al_8fddd1ab),
    .b(al_a7b01c14[2]),
    .c(al_df5cc0b8),
    .d(al_85a2bdb0[17]),
    .o(al_704d20e3[17]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(~D*~A)))"),
    .INIT(16'h0313))
    al_e0b21604 (
    .a(al_479534eb),
    .b(al_56afc96e),
    .c(al_28a777ae),
    .d(al_bdf9a7dd),
    .o(al_704d20e3[18]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    .INIT(16'hfbc8))
    al_4b3d3bd3 (
    .a(al_f7e849b8),
    .b(al_a7b01c14[2]),
    .c(al_2978bc8a),
    .d(al_85a2bdb0[20]),
    .o(al_704d20e3[20]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    .INIT(16'hfbc8))
    al_bdd7c8c2 (
    .a(al_b0c44f4),
    .b(al_a7b01c14[2]),
    .c(al_da3cc173),
    .d(al_85a2bdb0[21]),
    .o(al_704d20e3[21]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(~D*~A)))"),
    .INIT(16'h0313))
    al_86f7abae (
    .a(al_1bae5100),
    .b(al_8bc7d472),
    .c(al_55994c98),
    .d(al_bdf9a7dd),
    .o(al_704d20e3[22]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(~D*~A)))"),
    .INIT(16'h0313))
    al_30b1f9af (
    .a(al_c51bf9b),
    .b(al_136ceed1),
    .c(al_ffe7e6d4),
    .d(al_bdf9a7dd),
    .o(al_704d20e3[23]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_bc616bf5 (
    .a(al_f1e867e0),
    .b(al_a7b01c14[2]),
    .c(al_85a2bdb0[24]),
    .o(al_704d20e3[24]));
  AL_MAP_LUT6 #(
    .EQN("(~A*(B*~(C)*~(D)*~(E)*~(F)+B*C*~(D)*~(E)*~(F)+~(B)*~(C)*~(D)*E*~(F)+B*~(C)*~(D)*E*~(F)+~(B)*C*~(D)*E*~(F)+B*C*~(D)*E*~(F)+~(B)*~(C)*D*E*~(F)+B*~(C)*D*E*~(F)+~(B)*C*D*E*~(F)+B*C*D*E*~(F)+B*~(C)*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*~(C)*D*~(E)*F+B*~(C)*D*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*~(D)*E*F+B*~(C)*~(D)*E*F+B*C*~(D)*E*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'h5545554455550044))
    al_980c0369 (
    .a(al_1a551855),
    .b(al_de0f70d9),
    .c(al_8bea08a7),
    .d(al_85a2bdb0[3]),
    .e(al_85a2bdb0[4]),
    .f(al_85a2bdb0[6]),
    .o(al_170fdda));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7d9635f6 (
    .a(al_1ca0e00e),
    .b(al_c0a7a5f),
    .o(al_5493f072));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fffb3ba4 (
    .a(al_1edb758f[0]),
    .b(al_1edb758f[1]),
    .o(al_628a9731));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_e7655ee3 (
    .a(al_a2426a1),
    .b(al_cdace779),
    .c(al_24641d37),
    .d(al_501dbbdf),
    .o(al_b4eb77a8));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_252f1878 (
    .a(al_5493f072),
    .b(al_85a2bdb0[18]),
    .c(al_85a2bdb0[19]),
    .d(al_36a894af[10]),
    .e(al_36a894af[11]),
    .o(al_21c33d70));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_c1bf6fcf (
    .a(al_85a2bdb0[15]),
    .b(al_85a2bdb0[16]),
    .c(al_85a2bdb0[17]),
    .d(al_36a894af[7]),
    .e(al_36a894af[8]),
    .f(al_36a894af[9]),
    .o(al_ea118cf6));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    al_cf2ab1e (
    .a(al_b4eb77a8),
    .b(al_21c33d70),
    .c(al_ea118cf6),
    .o(al_71c814f5));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_26b5a4a4 (
    .a(al_6a6a2b33[1]),
    .b(al_6a6a2b33[3]),
    .c(al_6a6a2b33[4]),
    .d(al_85a2bdb0[16]),
    .e(al_85a2bdb0[18]),
    .f(al_85a2bdb0[19]),
    .o(al_a478b55f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_1fee1d9f (
    .a(al_501dbbdf),
    .b(al_bfc96350[0]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[0]),
    .f(al_d1fb6e0a[31]),
    .o(al_192eeeac[0]));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(F@D)*~(E@C))"),
    .INIT(64'h8000080000800008))
    al_8f3b330a (
    .a(al_a478b55f),
    .b(al_b3a31b1c),
    .c(al_6a6a2b33[0]),
    .d(al_6a6a2b33[2]),
    .e(al_85a2bdb0[15]),
    .f(al_85a2bdb0[17]),
    .o(al_d1df0873));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8116ea6c (
    .a(al_71c814f5),
    .b(al_b4eb77a8),
    .c(al_d1df0873),
    .o(al_e7747da7));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_ccd7d61b (
    .a(al_a62203af),
    .b(al_ebace85),
    .c(al_44595135),
    .d(al_523cde28),
    .o(al_4ed9ad89));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfac))
    al_26a14496 (
    .a(al_eebab250),
    .b(dBusAhb_HADDR[0]),
    .c(al_1edb758f[0]),
    .d(al_1edb758f[1]),
    .o(al_e3773112));
  AL_MAP_LUT5 #(
    .EQN("(C*(A*~(B)*~(D)*~(E)+~(A)*B*~(D)*~(E)+A*~(B)*D*~(E)+~(A)*~(B)*~(D)*E+A*~(B)*~(D)*E+A*B*~(D)*E+A*~(B)*D*E+~(A)*B*D*E))"),
    .INIT(32'h60b02060))
    al_17cc0087 (
    .a(al_f2330f79[0]),
    .b(al_18077581[0]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_de44ed56));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*A)*~(B)*~(D)+~(~C*A)*B*~(D)+~(~(~C*A))*B*D+~(~C*A)*B*D)"),
    .INIT(16'h330a))
    al_ecbf929b (
    .a(al_e3773112),
    .b(al_c0855656),
    .c(al_de44ed56),
    .d(al_b211b12d),
    .o(al_8221e5ce[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h02138a9b4657cedf))
    al_2c33870a (
    .a(al_e7747da7),
    .b(al_71c814f5),
    .c(al_8aeaa5c1[0]),
    .d(al_6fd79ca[0]),
    .e(al_4fd032af[0]),
    .f(al_81a1940d[0]),
    .o(al_18153c5c));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_fdd8a5b9 (
    .a(al_192eeeac[0]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[0]),
    .o(al_8aeaa5c1[0]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_9169780b (
    .a(al_18153c5c),
    .b(al_8221e5ce[0]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_7fc773bc (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .c(al_24ce3017[0]),
    .d(al_24ce3017[8]),
    .e(al_24ce3017[16]),
    .f(al_24ce3017[24]),
    .o(al_89494e6b));
  AL_MAP_LUT5 #(
    .EQN("(E*(B*~((~D*~C))*~(A)+B*(~D*~C)*~(A)+~(B)*(~D*~C)*A+B*(~D*~C)*A))"),
    .INIT(32'h444e0000))
    al_232e753f (
    .a(al_41e75372),
    .b(al_2af4b91),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_c0a7a5f),
    .o(al_781ea417));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_433870a2 (
    .a(al_41e75372),
    .b(al_c0a7a5f),
    .o(al_a559a13b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_798f3484 (
    .a(al_89494e6b),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[0]),
    .e(al_8900fb4e[0]),
    .f(al_d7ecfd18[0]),
    .o(al_6fd79ca[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_6dd725f2 (
    .a(al_501dbbdf),
    .b(al_bfc96350[10]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[10]),
    .f(al_d1fb6e0a[21]),
    .o(al_192eeeac[10]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_fe680007 (
    .a(al_e8e20039),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[10]),
    .o(al_bbc99cd7[10]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_55ca02ea (
    .a(al_192eeeac[10]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[10]),
    .o(al_8aeaa5c1[10]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~(~D*~C)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))"),
    .INIT(64'h0005111544455555))
    al_8406d862 (
    .a(al_68b1ca17),
    .b(al_5f3d7b85),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_24ce3017[10]),
    .f(al_24ce3017[26]),
    .o(al_d5e15803));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_a1b8c616 (
    .a(al_d5e15803),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[10]),
    .e(al_8900fb4e[10]),
    .f(al_d7ecfd18[10]),
    .o(al_6fd79ca[10]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_123841f6 (
    .a(al_f2330f79[10]),
    .b(al_18077581[10]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_fbf0401d));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_85496b45 (
    .a(al_fbf0401d),
    .b(dBusAhb_HADDR[10]),
    .c(al_354f5999),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[10]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010ba1ab515bf1fb))
    al_6ca1b862 (
    .a(al_e7747da7),
    .b(al_6fd79ca[10]),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[10]),
    .e(al_4fd032af[10]),
    .f(al_81a1940d[10]),
    .o(al_e8e20039));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_aa8baaab (
    .a(al_501dbbdf),
    .b(al_bfc96350[11]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[11]),
    .f(al_d1fb6e0a[20]),
    .o(al_192eeeac[11]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_36a87ee2 (
    .a(al_d2548651),
    .b(al_8221e5ce[11]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[11]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_5d78366d (
    .a(al_192eeeac[11]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[11]),
    .o(al_8aeaa5c1[11]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~(~D*~C)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))"),
    .INIT(64'h0005111544455555))
    al_9f00ce4d (
    .a(al_68b1ca17),
    .b(al_5f3d7b85),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_24ce3017[11]),
    .f(al_24ce3017[27]),
    .o(al_177c2401));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_7bf02eb7 (
    .a(al_177c2401),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[11]),
    .e(al_8900fb4e[11]),
    .f(al_d7ecfd18[11]),
    .o(al_6fd79ca[11]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_180ae080 (
    .a(al_f2330f79[11]),
    .b(al_18077581[11]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_bd6aed53));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_2d6cb6c4 (
    .a(al_5f34afe1),
    .b(al_bd6aed53),
    .c(dBusAhb_HADDR[11]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010ba1ab515bf1fb))
    al_7e2ed01a (
    .a(al_e7747da7),
    .b(al_6fd79ca[11]),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[11]),
    .e(al_4fd032af[11]),
    .f(al_81a1940d[11]),
    .o(al_d2548651));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_c7d20fc5 (
    .a(al_501dbbdf),
    .b(al_bfc96350[12]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[12]),
    .f(al_d1fb6e0a[19]),
    .o(al_192eeeac[12]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_3f569dca (
    .a(al_59035248),
    .b(al_8221e5ce[12]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[12]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_ac779f1d (
    .a(al_192eeeac[12]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[12]),
    .o(al_8aeaa5c1[12]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~(~D*~C)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))"),
    .INIT(64'h0005111544455555))
    al_bfbb9527 (
    .a(al_68b1ca17),
    .b(al_5f3d7b85),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_24ce3017[12]),
    .f(al_24ce3017[28]),
    .o(al_162afaa8));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_f46ce4d0 (
    .a(al_162afaa8),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[12]),
    .e(al_8900fb4e[12]),
    .f(al_d7ecfd18[12]),
    .o(al_6fd79ca[12]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_e3f33604 (
    .a(al_f2330f79[12]),
    .b(al_18077581[12]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_ba428019));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_98e7c7d4 (
    .a(al_63c14fc),
    .b(al_ba428019),
    .c(dBusAhb_HADDR[12]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010ba1ab515bf1fb))
    al_226e5746 (
    .a(al_e7747da7),
    .b(al_6fd79ca[12]),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[12]),
    .e(al_4fd032af[12]),
    .f(al_81a1940d[12]),
    .o(al_59035248));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_cee517c0 (
    .a(al_501dbbdf),
    .b(al_bfc96350[13]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[13]),
    .f(al_d1fb6e0a[18]),
    .o(al_192eeeac[13]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_6beba76 (
    .a(al_43aa4702),
    .b(al_8221e5ce[13]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[13]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_2c4132f9 (
    .a(al_192eeeac[13]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[13]),
    .o(al_8aeaa5c1[13]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~(~D*~C)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))"),
    .INIT(64'h0005111544455555))
    al_a198132b (
    .a(al_68b1ca17),
    .b(al_5f3d7b85),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_24ce3017[13]),
    .f(al_24ce3017[29]),
    .o(al_cae48ea4));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_fe5c5ada (
    .a(al_cae48ea4),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[13]),
    .e(al_8900fb4e[13]),
    .f(al_d7ecfd18[13]),
    .o(al_6fd79ca[13]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_fcbcb9f0 (
    .a(al_f2330f79[13]),
    .b(al_18077581[13]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_82238017));
  AL_MAP_LUT6 #(
    .EQN("~((~B*~(C*~(F@E)))*~(A)*~(D)+(~B*~(C*~(F@E)))*A*~(D)+~((~B*~(C*~(F@E))))*A*D+(~B*~(C*~(F@E)))*A*D)"),
    .INIT(64'h55fc55cc55cc55fc))
    al_9f8d19c9 (
    .a(al_85bef49),
    .b(al_82238017),
    .c(dBusAhb_HADDR[13]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010ba1ab515bf1fb))
    al_1c62e2d9 (
    .a(al_e7747da7),
    .b(al_6fd79ca[13]),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[13]),
    .e(al_4fd032af[13]),
    .f(al_81a1940d[13]),
    .o(al_43aa4702));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_f3298c2e (
    .a(al_501dbbdf),
    .b(al_bfc96350[14]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[14]),
    .f(al_d1fb6e0a[17]),
    .o(al_192eeeac[14]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_3bbc9289 (
    .a(al_b184fe5a),
    .b(al_8221e5ce[14]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[14]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_939446f6 (
    .a(al_192eeeac[14]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[14]),
    .o(al_8aeaa5c1[14]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~(~D*~C)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))"),
    .INIT(64'h0005111544455555))
    al_b9c7b603 (
    .a(al_68b1ca17),
    .b(al_5f3d7b85),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_24ce3017[14]),
    .f(al_24ce3017[30]),
    .o(al_cae74074));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_6c399c64 (
    .a(al_cae74074),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[14]),
    .e(al_8900fb4e[14]),
    .f(al_d7ecfd18[14]),
    .o(al_6fd79ca[14]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_127a8120 (
    .a(al_f2330f79[14]),
    .b(al_18077581[14]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_1a1782f2));
  AL_MAP_LUT6 #(
    .EQN("~((~B*~(C*~(F@E)))*~(A)*~(D)+(~B*~(C*~(F@E)))*A*~(D)+~((~B*~(C*~(F@E))))*A*D+(~B*~(C*~(F@E)))*A*D)"),
    .INIT(64'h55fc55cc55cc55fc))
    al_3c9e78ba (
    .a(al_94f9539),
    .b(al_1a1782f2),
    .c(dBusAhb_HADDR[14]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010ba1ab515bf1fb))
    al_d24b292e (
    .a(al_e7747da7),
    .b(al_6fd79ca[14]),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[14]),
    .e(al_4fd032af[14]),
    .f(al_81a1940d[14]),
    .o(al_b184fe5a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_44ba236e (
    .a(al_501dbbdf),
    .b(al_bfc96350[15]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[15]),
    .f(al_d1fb6e0a[16]),
    .o(al_192eeeac[15]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_6254a4c1 (
    .a(al_192eeeac[15]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[15]),
    .o(al_8aeaa5c1[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_62664166 (
    .a(al_286e2d87),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[15]),
    .e(al_8900fb4e[15]),
    .f(al_d7ecfd18[15]),
    .o(al_6fd79ca[15]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_a1839c29 (
    .a(al_f2330f79[15]),
    .b(al_18077581[15]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_a9bc0459));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_b716a1e7 (
    .a(al_a9bc0459),
    .b(dBusAhb_HADDR[15]),
    .c(al_f49386),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010ba1ab515bf1fb))
    al_682cfe98 (
    .a(al_e7747da7),
    .b(al_6fd79ca[15]),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[15]),
    .e(al_4fd032af[15]),
    .f(al_81a1940d[15]),
    .o(al_893ad164));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_a6ecc705 (
    .a(al_893ad164),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[15]),
    .o(al_bbc99cd7[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_57bbd94f (
    .a(al_501dbbdf),
    .b(al_bfc96350[16]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[15]),
    .f(al_d1fb6e0a[16]),
    .o(al_192eeeac[16]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_3a26391a (
    .a(al_e4ddc7f7),
    .b(al_8221e5ce[16]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[16]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_a28b5eff (
    .a(al_192eeeac[16]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[16]),
    .o(al_8aeaa5c1[16]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_f63c12d2 (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[16]),
    .e(al_8900fb4e[16]),
    .o(al_aa329d99));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_36fba8c6 (
    .a(al_aa329d99),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[16]),
    .e(al_d7ecfd18[16]),
    .o(al_6fd79ca[16]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_8f3e92c5 (
    .a(al_f2330f79[16]),
    .b(al_18077581[16]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_9d940ee8));
  AL_MAP_LUT6 #(
    .EQN("~((~B*~(C*~(F@E)))*~(A)*~(D)+(~B*~(C*~(F@E)))*A*~(D)+~((~B*~(C*~(F@E))))*A*D+(~B*~(C*~(F@E)))*A*D)"),
    .INIT(64'h55fc55cc55cc55fc))
    al_883f7d3d (
    .a(al_b44f8827),
    .b(al_9d940ee8),
    .c(dBusAhb_HADDR[16]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_3599ad7f (
    .a(al_6fd79ca[16]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[16]),
    .e(al_4fd032af[16]),
    .f(al_81a1940d[16]),
    .o(al_e4ddc7f7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_f581b56a (
    .a(al_501dbbdf),
    .b(al_bfc96350[17]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[14]),
    .f(al_d1fb6e0a[17]),
    .o(al_192eeeac[17]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_575d5a08 (
    .a(al_ad86ef7d),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[17]),
    .o(al_bbc99cd7[17]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_e9cd64d1 (
    .a(al_192eeeac[17]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[17]),
    .o(al_8aeaa5c1[17]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_fa205be (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[17]),
    .e(al_8900fb4e[17]),
    .o(al_45d4540c));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_1ec33384 (
    .a(al_45d4540c),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[17]),
    .e(al_d7ecfd18[17]),
    .o(al_6fd79ca[17]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_223a039d (
    .a(al_f2330f79[17]),
    .b(al_18077581[17]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_d71e234e));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_9d0b953 (
    .a(al_d71e234e),
    .b(dBusAhb_HADDR[17]),
    .c(al_daaf28b4),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_807e5759 (
    .a(al_6fd79ca[17]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[17]),
    .e(al_4fd032af[17]),
    .f(al_81a1940d[17]),
    .o(al_ad86ef7d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_bc7800c (
    .a(al_501dbbdf),
    .b(al_bfc96350[18]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[13]),
    .f(al_d1fb6e0a[18]),
    .o(al_192eeeac[18]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_8291cf38 (
    .a(al_aca053a7),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[18]),
    .o(al_bbc99cd7[18]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_1eb468c9 (
    .a(al_192eeeac[18]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[18]),
    .o(al_8aeaa5c1[18]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_46fc2b0a (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[18]),
    .e(al_8900fb4e[18]),
    .o(al_eb3feb88));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_9c4297bc (
    .a(al_eb3feb88),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[18]),
    .e(al_d7ecfd18[18]),
    .o(al_6fd79ca[18]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_a5916090 (
    .a(al_f2330f79[18]),
    .b(al_18077581[18]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_35e93aaa));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_5753aaed (
    .a(al_35e93aaa),
    .b(dBusAhb_HADDR[18]),
    .c(al_5c0f2717),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[18]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_b86d7d4e (
    .a(al_6fd79ca[18]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[18]),
    .e(al_4fd032af[18]),
    .f(al_81a1940d[18]),
    .o(al_aca053a7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_e1d64a2a (
    .a(al_501dbbdf),
    .b(al_bfc96350[19]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[12]),
    .f(al_d1fb6e0a[19]),
    .o(al_192eeeac[19]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_3395c6fb (
    .a(al_722a720c),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[19]),
    .o(al_bbc99cd7[19]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_47b2ce93 (
    .a(al_192eeeac[19]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[19]),
    .o(al_8aeaa5c1[19]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_d0f12014 (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[19]),
    .e(al_8900fb4e[19]),
    .o(al_7d5e05f7));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_7339134e (
    .a(al_7d5e05f7),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[19]),
    .e(al_d7ecfd18[19]),
    .o(al_6fd79ca[19]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_6cb1bdcc (
    .a(al_f2330f79[19]),
    .b(al_18077581[19]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_6b6f1ca9));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_cb0d1d54 (
    .a(al_6b6f1ca9),
    .b(dBusAhb_HADDR[19]),
    .c(al_8a79ceb4),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[19]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_822357dc (
    .a(al_6fd79ca[19]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[19]),
    .e(al_4fd032af[19]),
    .f(al_81a1940d[19]),
    .o(al_722a720c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_a383d746 (
    .a(al_501dbbdf),
    .b(al_bfc96350[1]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[1]),
    .f(al_d1fb6e0a[30]),
    .o(al_192eeeac[1]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_7890ae7d (
    .a(al_f41fca3f),
    .b(al_8221e5ce[1]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[1]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_ea698a5b (
    .a(al_192eeeac[1]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[1]),
    .o(al_8aeaa5c1[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_a200c0d0 (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .c(al_24ce3017[1]),
    .d(al_24ce3017[9]),
    .e(al_24ce3017[17]),
    .f(al_24ce3017[25]),
    .o(al_90b4cab0));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_b3910503 (
    .a(al_90b4cab0),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[1]),
    .e(al_8900fb4e[1]),
    .f(al_d7ecfd18[1]),
    .o(al_6fd79ca[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_cd9dc9d3 (
    .a(al_f2330f79[1]),
    .b(al_18077581[1]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_d83ea51));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_e01be907 (
    .a(al_f4418953),
    .b(al_d83ea51),
    .c(dBusAhb_HADDR[1]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h02138a9b4657cedf))
    al_2581ca38 (
    .a(al_e7747da7),
    .b(al_71c814f5),
    .c(al_8aeaa5c1[1]),
    .d(al_6fd79ca[1]),
    .e(al_4fd032af[1]),
    .f(al_81a1940d[1]),
    .o(al_f41fca3f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_a73661b1 (
    .a(al_501dbbdf),
    .b(al_bfc96350[20]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[11]),
    .f(al_d1fb6e0a[20]),
    .o(al_192eeeac[20]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_69d78f02 (
    .a(al_cdec8c3f),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[20]),
    .o(al_bbc99cd7[20]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_bec2307b (
    .a(al_192eeeac[20]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[20]),
    .o(al_8aeaa5c1[20]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_7131638c (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[20]),
    .e(al_8900fb4e[20]),
    .o(al_af9af7c7));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_eeaea769 (
    .a(al_af9af7c7),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[20]),
    .e(al_d7ecfd18[20]),
    .o(al_6fd79ca[20]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_456ffa6a (
    .a(al_f2330f79[20]),
    .b(al_18077581[20]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_94d4afd7));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_f5b447cc (
    .a(al_94d4afd7),
    .b(dBusAhb_HADDR[20]),
    .c(al_65a874f0),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[20]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_3ea5226 (
    .a(al_6fd79ca[20]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[20]),
    .e(al_4fd032af[20]),
    .f(al_81a1940d[20]),
    .o(al_cdec8c3f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_e1f5a309 (
    .a(al_501dbbdf),
    .b(al_bfc96350[21]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[10]),
    .f(al_d1fb6e0a[21]),
    .o(al_192eeeac[21]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_1e038eb4 (
    .a(al_c82d2f1e),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[21]),
    .o(al_bbc99cd7[21]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_79618381 (
    .a(al_192eeeac[21]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[21]),
    .o(al_8aeaa5c1[21]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_c2d110f0 (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[21]),
    .e(al_8900fb4e[21]),
    .o(al_2444302e));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_e2a9dfd9 (
    .a(al_2444302e),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[21]),
    .e(al_d7ecfd18[21]),
    .o(al_6fd79ca[21]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_815b79d6 (
    .a(al_f2330f79[21]),
    .b(al_18077581[21]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_8492fa3d));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_f5da022 (
    .a(al_8492fa3d),
    .b(dBusAhb_HADDR[21]),
    .c(al_80b925b7),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[21]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_4bbd54df (
    .a(al_6fd79ca[21]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[21]),
    .e(al_4fd032af[21]),
    .f(al_81a1940d[21]),
    .o(al_c82d2f1e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_360fb695 (
    .a(al_501dbbdf),
    .b(al_bfc96350[22]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[9]),
    .f(al_d1fb6e0a[22]),
    .o(al_192eeeac[22]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_119f0ea0 (
    .a(al_b67365e0),
    .b(al_8221e5ce[22]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[22]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_3755c483 (
    .a(al_192eeeac[22]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[22]),
    .o(al_8aeaa5c1[22]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_7d8a7d0f (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[22]),
    .e(al_8900fb4e[22]),
    .o(al_fa3c0cbe));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_fed90b53 (
    .a(al_fa3c0cbe),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[22]),
    .e(al_d7ecfd18[22]),
    .o(al_6fd79ca[22]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_eda17b48 (
    .a(al_f2330f79[22]),
    .b(al_18077581[22]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_13e3d996));
  AL_MAP_LUT6 #(
    .EQN("~((~B*~(C*~(F@E)))*~(A)*~(D)+(~B*~(C*~(F@E)))*A*~(D)+~((~B*~(C*~(F@E))))*A*D+(~B*~(C*~(F@E)))*A*D)"),
    .INIT(64'h55fc55cc55cc55fc))
    al_5119fee0 (
    .a(al_cb828215),
    .b(al_13e3d996),
    .c(dBusAhb_HADDR[22]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[22]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_b0822cc1 (
    .a(al_6fd79ca[22]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[22]),
    .e(al_4fd032af[22]),
    .f(al_81a1940d[22]),
    .o(al_b67365e0));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_d2b6c020 (
    .a(al_501dbbdf),
    .b(al_bfc96350[23]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[8]),
    .f(al_d1fb6e0a[23]),
    .o(al_192eeeac[23]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_198e9232 (
    .a(al_359eb4b6),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[23]),
    .o(al_bbc99cd7[23]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_cc709c4e (
    .a(al_192eeeac[23]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[23]),
    .o(al_8aeaa5c1[23]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_7d8203bb (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[23]),
    .e(al_8900fb4e[23]),
    .o(al_97c3f56c));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_ee3e0239 (
    .a(al_97c3f56c),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[23]),
    .e(al_d7ecfd18[23]),
    .o(al_6fd79ca[23]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_513feadb (
    .a(al_f2330f79[23]),
    .b(al_18077581[23]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_a3cc9c36));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_bdd91ce6 (
    .a(al_a3cc9c36),
    .b(dBusAhb_HADDR[23]),
    .c(al_ce80e68f),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[23]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_7fac4dd2 (
    .a(al_6fd79ca[23]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[23]),
    .e(al_4fd032af[23]),
    .f(al_81a1940d[23]),
    .o(al_359eb4b6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_e2a8e1d0 (
    .a(al_501dbbdf),
    .b(al_bfc96350[24]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[7]),
    .f(al_d1fb6e0a[24]),
    .o(al_192eeeac[24]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_7ddf629f (
    .a(al_b0f1a2c),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[24]),
    .o(al_bbc99cd7[24]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_d8536275 (
    .a(al_192eeeac[24]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[24]),
    .o(al_8aeaa5c1[24]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_9a8e886d (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[24]),
    .e(al_8900fb4e[24]),
    .o(al_ab419e9c));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_33a3abad (
    .a(al_ab419e9c),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[24]),
    .e(al_d7ecfd18[24]),
    .o(al_6fd79ca[24]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_c721ec41 (
    .a(al_f2330f79[24]),
    .b(al_18077581[24]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_4db2159c));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_13cb0aec (
    .a(al_4db2159c),
    .b(dBusAhb_HADDR[24]),
    .c(al_14816c03),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_de4442e4 (
    .a(al_6fd79ca[24]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[24]),
    .e(al_4fd032af[24]),
    .f(al_81a1940d[24]),
    .o(al_b0f1a2c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_278aaf9e (
    .a(al_501dbbdf),
    .b(al_bfc96350[25]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[6]),
    .f(al_d1fb6e0a[25]),
    .o(al_192eeeac[25]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_b51dbc19 (
    .a(al_1ae2d65b),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[25]),
    .o(al_bbc99cd7[25]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_31a325df (
    .a(al_192eeeac[25]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[25]),
    .o(al_8aeaa5c1[25]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_e2ce1664 (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[25]),
    .e(al_8900fb4e[25]),
    .o(al_deac45a7));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_6a314250 (
    .a(al_deac45a7),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[25]),
    .e(al_d7ecfd18[25]),
    .o(al_6fd79ca[25]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_88494028 (
    .a(al_f2330f79[25]),
    .b(al_18077581[25]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_819b6344));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_230aef56 (
    .a(al_819b6344),
    .b(dBusAhb_HADDR[25]),
    .c(al_6d174013),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_43fa10bb (
    .a(al_6fd79ca[25]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[25]),
    .e(al_4fd032af[25]),
    .f(al_81a1940d[25]),
    .o(al_1ae2d65b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_b248966 (
    .a(al_501dbbdf),
    .b(al_bfc96350[26]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[5]),
    .f(al_d1fb6e0a[26]),
    .o(al_192eeeac[26]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_dca118e3 (
    .a(al_2bed4baa),
    .b(al_8221e5ce[26]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[26]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_99062343 (
    .a(al_192eeeac[26]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[26]),
    .o(al_8aeaa5c1[26]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_5c34aaf7 (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[26]),
    .e(al_8900fb4e[26]),
    .o(al_73cede3c));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_9e9737cb (
    .a(al_73cede3c),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[26]),
    .e(al_d7ecfd18[26]),
    .o(al_6fd79ca[26]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_a28e711a (
    .a(al_f2330f79[26]),
    .b(al_18077581[26]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_4605c5c6));
  AL_MAP_LUT6 #(
    .EQN("~((~B*~(C*~(F@E)))*~(A)*~(D)+(~B*~(C*~(F@E)))*A*~(D)+~((~B*~(C*~(F@E))))*A*D+(~B*~(C*~(F@E)))*A*D)"),
    .INIT(64'h55fc55cc55cc55fc))
    al_7813ebd1 (
    .a(al_bb4f8966),
    .b(al_4605c5c6),
    .c(dBusAhb_HADDR[26]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_f0cff8de (
    .a(al_6fd79ca[26]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[26]),
    .e(al_4fd032af[26]),
    .f(al_81a1940d[26]),
    .o(al_2bed4baa));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_e2570f43 (
    .a(al_501dbbdf),
    .b(al_bfc96350[27]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[4]),
    .f(al_d1fb6e0a[27]),
    .o(al_192eeeac[27]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_23818b6 (
    .a(al_3813142e),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[27]),
    .o(al_bbc99cd7[27]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_dea0e34e (
    .a(al_192eeeac[27]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[27]),
    .o(al_8aeaa5c1[27]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_f823af1a (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[27]),
    .e(al_8900fb4e[27]),
    .o(al_362ab5dc));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_d9928480 (
    .a(al_362ab5dc),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[27]),
    .e(al_d7ecfd18[27]),
    .o(al_6fd79ca[27]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_755dedff (
    .a(al_f2330f79[27]),
    .b(al_18077581[27]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_b509771d));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_5418c086 (
    .a(al_b509771d),
    .b(dBusAhb_HADDR[27]),
    .c(al_70fea121),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_23045f23 (
    .a(al_6fd79ca[27]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[27]),
    .e(al_4fd032af[27]),
    .f(al_81a1940d[27]),
    .o(al_3813142e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_5eba5f3c (
    .a(al_501dbbdf),
    .b(al_bfc96350[28]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[3]),
    .f(al_d1fb6e0a[28]),
    .o(al_192eeeac[28]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_e808f515 (
    .a(al_cb20b6b1),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[28]),
    .o(al_bbc99cd7[28]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_a9bb8b4e (
    .a(al_192eeeac[28]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[28]),
    .o(al_8aeaa5c1[28]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_dc01b5d9 (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[28]),
    .e(al_8900fb4e[28]),
    .o(al_bfcbc23b));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_41dcab19 (
    .a(al_bfcbc23b),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[28]),
    .e(al_d7ecfd18[28]),
    .o(al_6fd79ca[28]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_5faef5 (
    .a(al_f2330f79[28]),
    .b(al_18077581[28]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_8e2aeac5));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_aaf2b176 (
    .a(al_8e2aeac5),
    .b(dBusAhb_HADDR[28]),
    .c(al_7750a3cd),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[28]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_dda41717 (
    .a(al_6fd79ca[28]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[28]),
    .e(al_4fd032af[28]),
    .f(al_81a1940d[28]),
    .o(al_cb20b6b1));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_51867694 (
    .a(al_501dbbdf),
    .b(al_bfc96350[29]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[2]),
    .f(al_d1fb6e0a[29]),
    .o(al_192eeeac[29]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_f6fed957 (
    .a(al_21fa7d09),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[29]),
    .o(al_bbc99cd7[29]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_7695faa1 (
    .a(al_192eeeac[29]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[29]),
    .o(al_8aeaa5c1[29]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_c1c69907 (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[29]),
    .e(al_8900fb4e[29]),
    .o(al_2beb9d89));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_9708bb42 (
    .a(al_2beb9d89),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[29]),
    .e(al_d7ecfd18[29]),
    .o(al_6fd79ca[29]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_6bf83a6b (
    .a(al_f2330f79[29]),
    .b(al_18077581[29]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_aae16022));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_93b6508f (
    .a(al_aae16022),
    .b(dBusAhb_HADDR[29]),
    .c(al_7b880725),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_ba223fea (
    .a(al_6fd79ca[29]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[29]),
    .e(al_4fd032af[29]),
    .f(al_81a1940d[29]),
    .o(al_21fa7d09));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_2c0aba8e (
    .a(al_501dbbdf),
    .b(al_bfc96350[2]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[2]),
    .f(al_d1fb6e0a[29]),
    .o(al_192eeeac[2]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_cddb3914 (
    .a(al_2e8a294f),
    .b(al_8221e5ce[2]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[2]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_39ebab34 (
    .a(al_192eeeac[2]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[2]),
    .o(al_8aeaa5c1[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_6d692378 (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .c(al_24ce3017[2]),
    .d(al_24ce3017[10]),
    .e(al_24ce3017[18]),
    .f(al_24ce3017[26]),
    .o(al_a7e3ba76));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_1612cc5e (
    .a(al_a7e3ba76),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[2]),
    .e(al_8900fb4e[2]),
    .f(al_d7ecfd18[2]),
    .o(al_6fd79ca[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_acefa81e (
    .a(al_f2330f79[2]),
    .b(al_18077581[2]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_93600cc2));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_57715968 (
    .a(al_a0c987d5),
    .b(al_93600cc2),
    .c(dBusAhb_HADDR[2]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h02138a9b4657cedf))
    al_63dc842b (
    .a(al_e7747da7),
    .b(al_71c814f5),
    .c(al_8aeaa5c1[2]),
    .d(al_6fd79ca[2]),
    .e(al_4fd032af[2]),
    .f(al_81a1940d[2]),
    .o(al_2e8a294f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_ae244404 (
    .a(al_501dbbdf),
    .b(al_bfc96350[30]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[1]),
    .f(al_d1fb6e0a[30]),
    .o(al_192eeeac[30]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_69294789 (
    .a(al_db9a596c),
    .b(al_8221e5ce[30]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[30]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_6666f760 (
    .a(al_192eeeac[30]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[30]),
    .o(al_8aeaa5c1[30]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_d0157797 (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[30]),
    .e(al_8900fb4e[30]),
    .o(al_5eff1a16));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_88237b02 (
    .a(al_5eff1a16),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[30]),
    .e(al_d7ecfd18[30]),
    .o(al_6fd79ca[30]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_390f0dbb (
    .a(al_f2330f79[30]),
    .b(al_18077581[30]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_a860806e));
  AL_MAP_LUT6 #(
    .EQN("~((~B*~(C*~(F@E)))*~(A)*~(D)+(~B*~(C*~(F@E)))*A*~(D)+~((~B*~(C*~(F@E))))*A*D+(~B*~(C*~(F@E)))*A*D)"),
    .INIT(64'h55fc55cc55cc55fc))
    al_556b3081 (
    .a(al_e9a9157c),
    .b(al_a860806e),
    .c(dBusAhb_HADDR[30]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_cdb17cea (
    .a(al_6fd79ca[30]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[30]),
    .e(al_4fd032af[30]),
    .f(al_81a1940d[30]),
    .o(al_db9a596c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeecee4c44ec444c))
    al_247fa8e1 (
    .a(al_501dbbdf),
    .b(al_bfc96350[31]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[0]),
    .f(al_d1fb6e0a[31]),
    .o(al_192eeeac[31]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_719d559a (
    .a(al_36a894af[13]),
    .b(al_36a894af[14]),
    .c(al_286e2d87),
    .o(al_7b1d42ce));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~A*~(D*C)))*~(B)+~E*(~A*~(D*C))*~(B)+~(~E)*(~A*~(D*C))*B+~E*(~A*~(D*C))*B)"),
    .INIT(32'h04443777))
    al_b75dda9c (
    .a(al_7b1d42ce),
    .b(al_781ea417),
    .c(al_36a894af[13]),
    .d(al_24ce3017[31]),
    .e(al_8900fb4e[31]),
    .o(al_4bbe4f7c));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    al_ff05f452 (
    .a(al_4bbe4f7c),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[31]),
    .e(al_d7ecfd18[31]),
    .o(al_6fd79ca[31]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_bff8ab10 (
    .a(al_f2330f79[31]),
    .b(al_18077581[31]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_18cae8b9));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_791493da (
    .a(al_ed766401),
    .b(al_18cae8b9),
    .c(dBusAhb_HADDR[31]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010dc1cd313df1fd))
    al_af39a76d (
    .a(al_6fd79ca[31]),
    .b(al_e7747da7),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[31]),
    .e(al_4fd032af[31]),
    .f(al_81a1940d[31]),
    .o(al_edead58e));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_62affe10 (
    .a(al_edead58e),
    .b(al_8221e5ce[31]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[31]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_f24996ac (
    .a(al_192eeeac[31]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[31]),
    .o(al_8aeaa5c1[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_a50ac139 (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .c(al_24ce3017[7]),
    .d(al_24ce3017[15]),
    .e(al_24ce3017[23]),
    .f(al_24ce3017[31]),
    .o(al_9dba4e2f));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_e075be9e (
    .a(al_9dba4e2f),
    .b(al_36a894af[12]),
    .c(al_36a894af[13]),
    .d(al_36a894af[14]),
    .o(al_68b1ca17));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cf74dfd7 (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .o(al_5f3d7b85));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~(~D*~C)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))"),
    .INIT(64'h0005111544455555))
    al_5ebfdc98 (
    .a(al_68b1ca17),
    .b(al_5f3d7b85),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_24ce3017[15]),
    .f(al_24ce3017[31]),
    .o(al_286e2d87));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_8471c7c9 (
    .a(al_501dbbdf),
    .b(al_bfc96350[3]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[3]),
    .f(al_d1fb6e0a[28]),
    .o(al_192eeeac[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_4effbcac (
    .a(al_618e5cf5),
    .b(al_8221e5ce[3]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_6fabdb46 (
    .a(al_192eeeac[3]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[3]),
    .o(al_8aeaa5c1[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_16bccaa1 (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .c(al_24ce3017[3]),
    .d(al_24ce3017[11]),
    .e(al_24ce3017[19]),
    .f(al_24ce3017[27]),
    .o(al_12251cca));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_71902b69 (
    .a(al_12251cca),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[3]),
    .e(al_8900fb4e[3]),
    .f(al_d7ecfd18[3]),
    .o(al_6fd79ca[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_21412bb2 (
    .a(al_f2330f79[3]),
    .b(al_18077581[3]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_63e36edf));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_49573ed7 (
    .a(al_1d8052bb),
    .b(al_63e36edf),
    .c(dBusAhb_HADDR[3]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h02138a9b4657cedf))
    al_a7aa555 (
    .a(al_e7747da7),
    .b(al_71c814f5),
    .c(al_8aeaa5c1[3]),
    .d(al_6fd79ca[3]),
    .e(al_4fd032af[3]),
    .f(al_81a1940d[3]),
    .o(al_618e5cf5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_fa983430 (
    .a(al_501dbbdf),
    .b(al_bfc96350[4]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[4]),
    .f(al_d1fb6e0a[27]),
    .o(al_192eeeac[4]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_52d3e578 (
    .a(al_3829588f),
    .b(al_8221e5ce[4]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[4]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_2a0043ab (
    .a(al_192eeeac[4]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[4]),
    .o(al_8aeaa5c1[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_c07aba85 (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .c(al_24ce3017[4]),
    .d(al_24ce3017[12]),
    .e(al_24ce3017[20]),
    .f(al_24ce3017[28]),
    .o(al_ed7763f6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_1cad07b9 (
    .a(al_ed7763f6),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[4]),
    .e(al_8900fb4e[4]),
    .f(al_d7ecfd18[4]),
    .o(al_6fd79ca[4]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_5aec2852 (
    .a(al_f2330f79[4]),
    .b(al_18077581[4]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_1ab00333));
  AL_MAP_LUT6 #(
    .EQN("~((~B*~(C*~(F@E)))*~(A)*~(D)+(~B*~(C*~(F@E)))*A*~(D)+~((~B*~(C*~(F@E))))*A*D+(~B*~(C*~(F@E)))*A*D)"),
    .INIT(64'h55fc55cc55cc55fc))
    al_2ea4f332 (
    .a(al_e0306332),
    .b(al_1ab00333),
    .c(dBusAhb_HADDR[4]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h02138a9b4657cedf))
    al_68cd56d8 (
    .a(al_e7747da7),
    .b(al_71c814f5),
    .c(al_8aeaa5c1[4]),
    .d(al_6fd79ca[4]),
    .e(al_4fd032af[4]),
    .f(al_81a1940d[4]),
    .o(al_3829588f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_7dee673e (
    .a(al_501dbbdf),
    .b(al_bfc96350[5]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[5]),
    .f(al_d1fb6e0a[26]),
    .o(al_192eeeac[5]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_50b1356c (
    .a(al_90adbe55),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[5]),
    .o(al_bbc99cd7[5]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_ae7d9772 (
    .a(al_192eeeac[5]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[5]),
    .o(al_8aeaa5c1[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_aec7285f (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .c(al_24ce3017[5]),
    .d(al_24ce3017[13]),
    .e(al_24ce3017[21]),
    .f(al_24ce3017[29]),
    .o(al_2295e150));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_9281e502 (
    .a(al_2295e150),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[5]),
    .e(al_8900fb4e[5]),
    .f(al_d7ecfd18[5]),
    .o(al_6fd79ca[5]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_4bb049ca (
    .a(al_f2330f79[5]),
    .b(al_18077581[5]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_bef23915));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_3c4c2783 (
    .a(al_bef23915),
    .b(dBusAhb_HADDR[5]),
    .c(al_75b09ba0),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h02138a9b4657cedf))
    al_23445c2b (
    .a(al_e7747da7),
    .b(al_71c814f5),
    .c(al_8aeaa5c1[5]),
    .d(al_6fd79ca[5]),
    .e(al_4fd032af[5]),
    .f(al_81a1940d[5]),
    .o(al_90adbe55));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_3f944eb2 (
    .a(al_501dbbdf),
    .b(al_bfc96350[6]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[6]),
    .f(al_d1fb6e0a[25]),
    .o(al_192eeeac[6]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_aac3768 (
    .a(al_5278baaa),
    .b(al_8221e5ce[6]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[6]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_5d1aea76 (
    .a(al_192eeeac[6]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[6]),
    .o(al_8aeaa5c1[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_547af9de (
    .a(al_70c1ae82[0]),
    .b(al_70c1ae82[1]),
    .c(al_24ce3017[6]),
    .d(al_24ce3017[14]),
    .e(al_24ce3017[22]),
    .f(al_24ce3017[30]),
    .o(al_3386891f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_343ba60d (
    .a(al_3386891f),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[6]),
    .e(al_8900fb4e[6]),
    .f(al_d7ecfd18[6]),
    .o(al_6fd79ca[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_2c7dbdd9 (
    .a(al_f2330f79[6]),
    .b(al_18077581[6]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_495a58bd));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_951290ad (
    .a(al_bb5767ca),
    .b(al_495a58bd),
    .c(dBusAhb_HADDR[6]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h02138a9b4657cedf))
    al_ad8629fc (
    .a(al_e7747da7),
    .b(al_71c814f5),
    .c(al_8aeaa5c1[6]),
    .d(al_6fd79ca[6]),
    .e(al_4fd032af[6]),
    .f(al_81a1940d[6]),
    .o(al_5278baaa));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_33c4d930 (
    .a(al_501dbbdf),
    .b(al_bfc96350[7]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[7]),
    .f(al_d1fb6e0a[24]),
    .o(al_192eeeac[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_6a1b5bb6 (
    .a(al_192eeeac[7]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[7]),
    .o(al_8aeaa5c1[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_ca09c3b9 (
    .a(al_9dba4e2f),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[7]),
    .e(al_8900fb4e[7]),
    .f(al_d7ecfd18[7]),
    .o(al_6fd79ca[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_e7d89583 (
    .a(al_f2330f79[7]),
    .b(al_18077581[7]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_26f7099d));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_e29542b0 (
    .a(al_83268b9b),
    .b(al_26f7099d),
    .c(dBusAhb_HADDR[7]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h02138a9b4657cedf))
    al_377c8398 (
    .a(al_e7747da7),
    .b(al_71c814f5),
    .c(al_8aeaa5c1[7]),
    .d(al_6fd79ca[7]),
    .e(al_4fd032af[7]),
    .f(al_81a1940d[7]),
    .o(al_7a187fb8));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_ab3a09e7 (
    .a(al_7a187fb8),
    .b(al_8221e5ce[7]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_b04f6e02 (
    .a(al_501dbbdf),
    .b(al_bfc96350[8]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[8]),
    .f(al_d1fb6e0a[23]),
    .o(al_192eeeac[8]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_8bc1ad87 (
    .a(al_63f22050),
    .b(al_4ed9ad89),
    .c(al_8221e5ce[8]),
    .o(al_bbc99cd7[8]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_4f5d049d (
    .a(al_192eeeac[8]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[8]),
    .o(al_8aeaa5c1[8]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~(~D*~C)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))"),
    .INIT(64'h0005111544455555))
    al_2e8d4734 (
    .a(al_68b1ca17),
    .b(al_5f3d7b85),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_24ce3017[8]),
    .f(al_24ce3017[24]),
    .o(al_541e0d8b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_e167bdb2 (
    .a(al_541e0d8b),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[8]),
    .e(al_8900fb4e[8]),
    .f(al_d7ecfd18[8]),
    .o(al_6fd79ca[8]));
  AL_MAP_LUT5 #(
    .EQN("(C*(~(A)*~(B)*~(D)*~(E)+A*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+~(A)*B*D*~(E)+A*B*D*~(E)+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h9040d090))
    al_93bed8f9 (
    .a(al_f2330f79[8]),
    .b(al_18077581[8]),
    .c(al_628a9731),
    .d(al_bb6625de[0]),
    .e(al_bb6625de[1]),
    .o(al_b950f9ad));
  AL_MAP_LUT6 #(
    .EQN("~((~A*~(B*~(F@E)))*~(C)*~(D)+(~A*~(B*~(F@E)))*C*~(D)+~((~A*~(B*~(F@E))))*C*D+(~A*~(B*~(F@E)))*C*D)"),
    .INIT(64'h0fee0faa0faa0fee))
    al_d89c932c (
    .a(al_b950f9ad),
    .b(dBusAhb_HADDR[8]),
    .c(al_26af78f7),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010ba1ab515bf1fb))
    al_c353ba7a (
    .a(al_e7747da7),
    .b(al_6fd79ca[8]),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[8]),
    .e(al_4fd032af[8]),
    .f(al_81a1940d[8]),
    .o(al_63f22050));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'heeec44ecee4c444c))
    al_e4295eef (
    .a(al_501dbbdf),
    .b(al_bfc96350[9]),
    .c(al_727d2e98[0]),
    .d(al_727d2e98[1]),
    .e(al_d1fb6e0a[9]),
    .f(al_d1fb6e0a[22]),
    .o(al_192eeeac[9]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_2157a2ef (
    .a(al_5bc78df0),
    .b(al_8221e5ce[9]),
    .c(al_4ed9ad89),
    .o(al_bbc99cd7[9]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((C*B))+A*D*~((C*B))+~(A)*D*(C*B)+A*D*(C*B))"),
    .INIT(16'hea2a))
    al_59977ed9 (
    .a(al_192eeeac[9]),
    .b(al_b2739b77),
    .c(al_501dbbdf),
    .d(al_ec26021c[9]),
    .o(al_8aeaa5c1[9]));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~(~D*~C)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))"),
    .INIT(64'h0005111544455555))
    al_c4bb931a (
    .a(al_68b1ca17),
    .b(al_5f3d7b85),
    .c(al_36a894af[12]),
    .d(al_36a894af[13]),
    .e(al_24ce3017[9]),
    .f(al_24ce3017[25]),
    .o(al_692e1afb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf737f434c707c404))
    al_4c96fc32 (
    .a(al_692e1afb),
    .b(al_781ea417),
    .c(al_a559a13b),
    .d(al_71c7f8f0[9]),
    .e(al_8900fb4e[9]),
    .f(al_d7ecfd18[9]),
    .o(al_6fd79ca[9]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*B*C*D)"),
    .INIT(16'h94d9))
    al_e9d3e6f2 (
    .a(al_f2330f79[9]),
    .b(al_18077581[9]),
    .c(al_bb6625de[0]),
    .d(al_bb6625de[1]),
    .o(al_972ccb4f));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*~(A)*~(D)+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*~(D)+~(~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F))*A*D+~(~(B)*C*~(E)*~(F)+B*C*~(E)*~(F)+B*~(C)*~(E)*F+B*C*~(E)*F+~(B)*C*E*F+B*C*E*F)*A*D)"),
    .INIT(64'h55f055cc550055f0))
    al_e74df9d6 (
    .a(al_29a1a38f),
    .b(al_972ccb4f),
    .c(dBusAhb_HADDR[9]),
    .d(al_b211b12d),
    .e(al_1edb758f[0]),
    .f(al_1edb758f[1]),
    .o(al_8221e5ce[9]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h010ba1ab515bf1fb))
    al_12ddcd3d (
    .a(al_e7747da7),
    .b(al_6fd79ca[9]),
    .c(al_71c814f5),
    .d(al_8aeaa5c1[9]),
    .e(al_4fd032af[9]),
    .f(al_81a1940d[9]),
    .o(al_5bc78df0));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_9cc1d17 (
    .a(al_5493f072),
    .b(al_85a2bdb0[23]),
    .c(al_85a2bdb0[24]),
    .d(al_36a894af[10]),
    .e(al_36a894af[11]),
    .o(al_b669e5e6));
  AL_MAP_LUT6 #(
    .EQN("~((F*E*D*B)*~(C)*~(A)+(F*E*D*B)*C*~(A)+~((F*E*D*B))*C*A+(F*E*D*B)*C*A)"),
    .INIT(64'h1b5f5f5f5f5f5f5f))
    al_a901001b (
    .a(al_e8448fdd),
    .b(al_df2df2f9),
    .c(al_1b14c7a0),
    .d(al_cdace779),
    .e(al_24641d37),
    .f(al_501dbbdf),
    .o(al_467f9b5e));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_d2e23c0 (
    .a(al_358f5bea),
    .b(al_ebace85),
    .c(al_44595135),
    .d(al_523cde28),
    .o(al_fc39fece));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_7ff7a982 (
    .a(al_467f9b5e),
    .b(al_e8448fdd),
    .c(al_8aeaa5c1[0]),
    .d(al_6fd79ca[0]),
    .e(al_4fd032af[0]),
    .f(al_fe073fc9[0]),
    .o(al_f48cb7f2));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_9613f729 (
    .a(al_f48cb7f2),
    .b(al_8221e5ce[0]),
    .c(al_fc39fece),
    .o(al_52ea52d7[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_cb4771d2 (
    .a(al_85a2bdb0[20]),
    .b(al_85a2bdb0[21]),
    .c(al_85a2bdb0[22]),
    .d(al_36a894af[7]),
    .e(al_36a894af[8]),
    .f(al_36a894af[9]),
    .o(al_a8b9ff36));
  AL_MAP_LUT6 #(
    .EQN("(~(C*B)*~(F*E*D*A))"),
    .INIT(64'h153f3f3f3f3f3f3f))
    al_4f570200 (
    .a(al_df2df2f9),
    .b(al_b669e5e6),
    .c(al_a8b9ff36),
    .d(al_cdace779),
    .e(al_24641d37),
    .f(al_501dbbdf),
    .o(al_e8448fdd));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_396f6fa1 (
    .a(al_6a6a2b33[1]),
    .b(al_6a6a2b33[3]),
    .c(al_6a6a2b33[4]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[23]),
    .f(al_85a2bdb0[24]),
    .o(al_71cdacfd));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(F@D)*~(E@C))"),
    .INIT(64'h8000080000800008))
    al_4e508e6f (
    .a(al_71cdacfd),
    .b(al_b3a31b1c),
    .c(al_6a6a2b33[0]),
    .d(al_6a6a2b33[2]),
    .e(al_85a2bdb0[20]),
    .f(al_85a2bdb0[22]),
    .o(al_1b14c7a0));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_df999dac (
    .a(al_6fd79ca[10]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[10]),
    .e(al_4fd032af[10]),
    .f(al_fe073fc9[10]),
    .o(al_12004dbe));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_3b360bc0 (
    .a(al_12004dbe),
    .b(al_fc39fece),
    .c(al_8221e5ce[10]),
    .o(al_52ea52d7[10]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_b4f12991 (
    .a(al_6fd79ca[11]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[11]),
    .e(al_4fd032af[11]),
    .f(al_fe073fc9[11]),
    .o(al_f7851a1a));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_d984020a (
    .a(al_f7851a1a),
    .b(al_8221e5ce[11]),
    .c(al_fc39fece),
    .o(al_52ea52d7[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_c2e2dfe8 (
    .a(al_6fd79ca[12]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[12]),
    .e(al_4fd032af[12]),
    .f(al_fe073fc9[12]),
    .o(al_d6db317));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_de96ee30 (
    .a(al_d6db317),
    .b(al_8221e5ce[12]),
    .c(al_fc39fece),
    .o(al_52ea52d7[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_9fe84ca6 (
    .a(al_6fd79ca[13]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[13]),
    .e(al_4fd032af[13]),
    .f(al_fe073fc9[13]),
    .o(al_d2b99696));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_3b231fc2 (
    .a(al_d2b99696),
    .b(al_8221e5ce[13]),
    .c(al_fc39fece),
    .o(al_52ea52d7[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_546753f5 (
    .a(al_6fd79ca[14]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[14]),
    .e(al_4fd032af[14]),
    .f(al_fe073fc9[14]),
    .o(al_477e72e5));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_d0a9e17a (
    .a(al_477e72e5),
    .b(al_8221e5ce[14]),
    .c(al_fc39fece),
    .o(al_52ea52d7[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_c805eb3a (
    .a(al_6fd79ca[15]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[15]),
    .e(al_4fd032af[15]),
    .f(al_fe073fc9[15]),
    .o(al_25614342));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_d97e943c (
    .a(al_25614342),
    .b(al_fc39fece),
    .c(al_8221e5ce[15]),
    .o(al_52ea52d7[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_518a72e0 (
    .a(al_6fd79ca[16]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[16]),
    .e(al_4fd032af[16]),
    .f(al_fe073fc9[16]),
    .o(al_9328cdb4));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_7af88c75 (
    .a(al_9328cdb4),
    .b(al_8221e5ce[16]),
    .c(al_fc39fece),
    .o(al_52ea52d7[16]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_93183fb2 (
    .a(al_6fd79ca[17]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[17]),
    .e(al_4fd032af[17]),
    .f(al_fe073fc9[17]),
    .o(al_3e17171c));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_7be2cc54 (
    .a(al_3e17171c),
    .b(al_fc39fece),
    .c(al_8221e5ce[17]),
    .o(al_52ea52d7[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_8b37ff12 (
    .a(al_6fd79ca[18]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[18]),
    .e(al_4fd032af[18]),
    .f(al_fe073fc9[18]),
    .o(al_1dab850a));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_324a819a (
    .a(al_1dab850a),
    .b(al_fc39fece),
    .c(al_8221e5ce[18]),
    .o(al_52ea52d7[18]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_d050aeeb (
    .a(al_6fd79ca[19]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[19]),
    .e(al_4fd032af[19]),
    .f(al_fe073fc9[19]),
    .o(al_cbe76bf6));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_b9dafa6e (
    .a(al_cbe76bf6),
    .b(al_fc39fece),
    .c(al_8221e5ce[19]),
    .o(al_52ea52d7[19]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_c291bc7a (
    .a(al_467f9b5e),
    .b(al_e8448fdd),
    .c(al_8aeaa5c1[1]),
    .d(al_6fd79ca[1]),
    .e(al_4fd032af[1]),
    .f(al_fe073fc9[1]),
    .o(al_81feda1d));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_b075f343 (
    .a(al_81feda1d),
    .b(al_8221e5ce[1]),
    .c(al_fc39fece),
    .o(al_52ea52d7[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_54fadb44 (
    .a(al_6fd79ca[20]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[20]),
    .e(al_4fd032af[20]),
    .f(al_fe073fc9[20]),
    .o(al_e3e05361));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_91f96450 (
    .a(al_e3e05361),
    .b(al_fc39fece),
    .c(al_8221e5ce[20]),
    .o(al_52ea52d7[20]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_bc541ece (
    .a(al_6fd79ca[21]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[21]),
    .e(al_4fd032af[21]),
    .f(al_fe073fc9[21]),
    .o(al_bee19057));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_4d53a1f2 (
    .a(al_bee19057),
    .b(al_fc39fece),
    .c(al_8221e5ce[21]),
    .o(al_52ea52d7[21]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_4c7d727c (
    .a(al_6fd79ca[22]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[22]),
    .e(al_4fd032af[22]),
    .f(al_fe073fc9[22]),
    .o(al_f176a1bb));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_229925a5 (
    .a(al_f176a1bb),
    .b(al_8221e5ce[22]),
    .c(al_fc39fece),
    .o(al_52ea52d7[22]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_2a70feba (
    .a(al_6fd79ca[23]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[23]),
    .e(al_4fd032af[23]),
    .f(al_fe073fc9[23]),
    .o(al_7989383a));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_e02c4530 (
    .a(al_7989383a),
    .b(al_fc39fece),
    .c(al_8221e5ce[23]),
    .o(al_52ea52d7[23]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_1bd5c29a (
    .a(al_6fd79ca[24]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[24]),
    .e(al_4fd032af[24]),
    .f(al_fe073fc9[24]),
    .o(al_36f32db5));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_facc09da (
    .a(al_36f32db5),
    .b(al_fc39fece),
    .c(al_8221e5ce[24]),
    .o(al_52ea52d7[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_9710d747 (
    .a(al_6fd79ca[25]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[25]),
    .e(al_4fd032af[25]),
    .f(al_fe073fc9[25]),
    .o(al_dea79dda));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_48872f5b (
    .a(al_dea79dda),
    .b(al_fc39fece),
    .c(al_8221e5ce[25]),
    .o(al_52ea52d7[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_5f9af51b (
    .a(al_6fd79ca[26]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[26]),
    .e(al_4fd032af[26]),
    .f(al_fe073fc9[26]),
    .o(al_74b0792c));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_5b8c5e86 (
    .a(al_74b0792c),
    .b(al_8221e5ce[26]),
    .c(al_fc39fece),
    .o(al_52ea52d7[26]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_d6446abe (
    .a(al_6fd79ca[27]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[27]),
    .e(al_4fd032af[27]),
    .f(al_fe073fc9[27]),
    .o(al_88c7c32a));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_8cf484ae (
    .a(al_88c7c32a),
    .b(al_fc39fece),
    .c(al_8221e5ce[27]),
    .o(al_52ea52d7[27]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_ef2795c5 (
    .a(al_6fd79ca[28]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[28]),
    .e(al_4fd032af[28]),
    .f(al_fe073fc9[28]),
    .o(al_d358a549));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_237c3061 (
    .a(al_d358a549),
    .b(al_fc39fece),
    .c(al_8221e5ce[28]),
    .o(al_52ea52d7[28]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_d2854ff0 (
    .a(al_6fd79ca[29]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[29]),
    .e(al_4fd032af[29]),
    .f(al_fe073fc9[29]),
    .o(al_16eb3ffd));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_9a606b2b (
    .a(al_16eb3ffd),
    .b(al_fc39fece),
    .c(al_8221e5ce[29]),
    .o(al_52ea52d7[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_bd92521b (
    .a(al_467f9b5e),
    .b(al_e8448fdd),
    .c(al_8aeaa5c1[2]),
    .d(al_6fd79ca[2]),
    .e(al_4fd032af[2]),
    .f(al_fe073fc9[2]),
    .o(al_433e30e8));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_f0b47126 (
    .a(al_433e30e8),
    .b(al_8221e5ce[2]),
    .c(al_fc39fece),
    .o(al_52ea52d7[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_1f0761e3 (
    .a(al_6fd79ca[30]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[30]),
    .e(al_4fd032af[30]),
    .f(al_fe073fc9[30]),
    .o(al_95046a85));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_694a5648 (
    .a(al_95046a85),
    .b(al_8221e5ce[30]),
    .c(al_fc39fece),
    .o(al_52ea52d7[30]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_5beb41ca (
    .a(al_6fd79ca[31]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[31]),
    .e(al_4fd032af[31]),
    .f(al_fe073fc9[31]),
    .o(al_89d8e10c));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_b2b563c5 (
    .a(al_89d8e10c),
    .b(al_8221e5ce[31]),
    .c(al_fc39fece),
    .o(al_52ea52d7[31]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_54ab0212 (
    .a(al_467f9b5e),
    .b(al_e8448fdd),
    .c(al_8aeaa5c1[3]),
    .d(al_6fd79ca[3]),
    .e(al_4fd032af[3]),
    .f(al_fe073fc9[3]),
    .o(al_51a7aab3));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_be2e45eb (
    .a(al_51a7aab3),
    .b(al_8221e5ce[3]),
    .c(al_fc39fece),
    .o(al_52ea52d7[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_34891f2e (
    .a(al_467f9b5e),
    .b(al_e8448fdd),
    .c(al_8aeaa5c1[4]),
    .d(al_6fd79ca[4]),
    .e(al_4fd032af[4]),
    .f(al_fe073fc9[4]),
    .o(al_1a113696));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_f7f032af (
    .a(al_1a113696),
    .b(al_8221e5ce[4]),
    .c(al_fc39fece),
    .o(al_52ea52d7[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_4e853e4d (
    .a(al_467f9b5e),
    .b(al_e8448fdd),
    .c(al_8aeaa5c1[5]),
    .d(al_6fd79ca[5]),
    .e(al_4fd032af[5]),
    .f(al_fe073fc9[5]),
    .o(al_568ed982));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_2450f677 (
    .a(al_568ed982),
    .b(al_fc39fece),
    .c(al_8221e5ce[5]),
    .o(al_52ea52d7[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_f9dfb9f8 (
    .a(al_467f9b5e),
    .b(al_e8448fdd),
    .c(al_8aeaa5c1[6]),
    .d(al_6fd79ca[6]),
    .e(al_4fd032af[6]),
    .f(al_fe073fc9[6]),
    .o(al_53750577));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_d084b4de (
    .a(al_53750577),
    .b(al_8221e5ce[6]),
    .c(al_fc39fece),
    .o(al_52ea52d7[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_d2a5ae5a (
    .a(al_467f9b5e),
    .b(al_e8448fdd),
    .c(al_8aeaa5c1[7]),
    .d(al_6fd79ca[7]),
    .e(al_4fd032af[7]),
    .f(al_fe073fc9[7]),
    .o(al_79961e57));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_64a5fa08 (
    .a(al_79961e57),
    .b(al_8221e5ce[7]),
    .c(al_fc39fece),
    .o(al_52ea52d7[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_adeffb48 (
    .a(al_6fd79ca[8]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[8]),
    .e(al_4fd032af[8]),
    .f(al_fe073fc9[8]),
    .o(al_406777f2));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_96f84937 (
    .a(al_406777f2),
    .b(al_fc39fece),
    .c(al_8221e5ce[8]),
    .o(al_52ea52d7[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_1693f92c (
    .a(al_6fd79ca[9]),
    .b(al_467f9b5e),
    .c(al_e8448fdd),
    .d(al_8aeaa5c1[9]),
    .e(al_4fd032af[9]),
    .f(al_fe073fc9[9]),
    .o(al_7fc6feef));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    al_5e9978a8 (
    .a(al_7fc6feef),
    .b(al_8221e5ce[9]),
    .c(al_fc39fece),
    .o(al_52ea52d7[9]));
  AL_DFF_X al_7d56af15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c0c7b1b4),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebace85));
  AL_DFF_X al_2b42aeb6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_4a753b95[11]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b2d5c80));
  AL_DFF_X al_e6157e0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_566f1754),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6715e869));
  AL_DFF_X al_77e16d60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2434efda),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_39cb3b56));
  AL_DFF_X al_ef0786a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c4aa9af),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbdc72d2));
  AL_DFF_X al_797cb85e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bb2524be),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8bf5da64));
  AL_DFF_X al_e47a06a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_361dafb5),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5b8f9ea));
  AL_DFF_X al_d133e6ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_66fb6e33),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9a05e7eb));
  AL_DFF_X al_c26c4cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b63bb946),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e46fbe7));
  AL_DFF_X al_7439398d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_24a3e858),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bcd349b));
  AL_DFF_X al_d2af640a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c52295d9),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32fedef4));
  AL_DFF_X al_ad0bc4a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[5]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWRITE));
  AL_DFF_X al_d341b1bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_da9c21fb),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86fb87b9));
  AL_DFF_X al_7ed32b3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_170fdda),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44595135));
  AL_DFF_X al_eeab19e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b8ccdc1c),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36962d69));
  AL_DFF_X al_54f88abd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_192b30b5),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aded6184));
  AL_DFF_X al_638a90ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_118827bc),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_df7b4407));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_88c333f7 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[31]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_60dd36d7),
    .o(al_f2330f79[31]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_7cc62d66 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[22]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_ffc4fe26),
    .o(al_f2330f79[22]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_73ea55a9 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[21]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_658bb789),
    .o(al_f2330f79[21]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_fde33705 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[20]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_a831c176),
    .o(al_f2330f79[20]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_7ae2f7fd (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[19]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_c7df4b4d),
    .o(al_f2330f79[19]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_d93cb786 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[18]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_3b0f4da7),
    .o(al_f2330f79[18]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_d93ab7a3 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[17]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_d76255c5),
    .o(al_f2330f79[17]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_19433fc8 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[16]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_7d27d680),
    .o(al_f2330f79[16]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_8f566adc (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[15]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_f61ec828),
    .o(al_f2330f79[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_f7b3de40 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[14]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_7e6320f4),
    .o(al_f2330f79[14]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_5cde846 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[13]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_e6455839),
    .o(al_f2330f79[13]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_650d2641 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[30]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_f1bb92e9),
    .o(al_f2330f79[30]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_48feb2ce (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[12]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_d00a6f56),
    .o(al_f2330f79[12]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_3ac1c38a (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[11]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_3ebb68c3),
    .o(al_f2330f79[11]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_cdfb9931 (
    .a(al_e03b3126[30]),
    .b(al_9bf95cff[10]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_98804c07),
    .o(al_f2330f79[10]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_63939fda (
    .a(al_e03b3126[29]),
    .b(al_9bf95cff[9]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_6d92b3c6),
    .o(al_f2330f79[9]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_42a64dc4 (
    .a(al_e03b3126[28]),
    .b(al_9bf95cff[8]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_bdb28b76),
    .o(al_f2330f79[8]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_eda3e4f4 (
    .a(al_e03b3126[27]),
    .b(al_9bf95cff[7]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_73fb1ee5),
    .o(al_f2330f79[7]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_a56f5fe3 (
    .a(al_e03b3126[26]),
    .b(al_9bf95cff[6]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_33a2911e),
    .o(al_f2330f79[6]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_1c8ca252 (
    .a(al_e03b3126[25]),
    .b(al_9bf95cff[5]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_8a841cb4),
    .o(al_f2330f79[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f5533000f5533ff))
    al_e332b877 (
    .a(al_e03b3126[11]),
    .b(al_e03b3126[24]),
    .c(al_9bf95cff[4]),
    .d(al_a1e88c0c[0]),
    .e(al_a1e88c0c[1]),
    .f(al_c861c8f0),
    .o(al_f2330f79[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f5533000f5533ff))
    al_f28bfe2c (
    .a(al_e03b3126[10]),
    .b(al_e03b3126[23]),
    .c(al_9bf95cff[3]),
    .d(al_a1e88c0c[0]),
    .e(al_a1e88c0c[1]),
    .f(al_76a52f3d),
    .o(al_f2330f79[3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_15563e27 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[29]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_3626cb0),
    .o(al_f2330f79[29]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f5533000f5533ff))
    al_85bced8f (
    .a(al_e03b3126[9]),
    .b(al_e03b3126[22]),
    .c(al_9bf95cff[2]),
    .d(al_a1e88c0c[0]),
    .e(al_a1e88c0c[1]),
    .f(al_bf952132),
    .o(al_f2330f79[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0f5533000f5533ff))
    al_c3009a0a (
    .a(al_e03b3126[8]),
    .b(al_e03b3126[21]),
    .c(al_9bf95cff[1]),
    .d(al_a1e88c0c[0]),
    .e(al_a1e88c0c[1]),
    .f(al_2370214),
    .o(al_f2330f79[1]));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h2be8))
    al_341faa2 (
    .a(dBusAhb_HADDR[31]),
    .b(al_f2330f79[31]),
    .c(al_18077581[31]),
    .d(al_aded6184),
    .o(al_eebab250));
  AL_MAP_LUT6 #(
    .EQN("((D@C)*(F@B)*(E@A))"),
    .INIT(64'h0110022004400880))
    al_f1d062be (
    .a(al_f2330f79[3]),
    .b(al_f2330f79[0]),
    .c(al_f2330f79[25]),
    .d(al_18077581[25]),
    .e(al_18077581[3]),
    .f(al_18077581[0]),
    .o(al_e2608c20));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    al_6edecb1a (
    .a(al_f2330f79[31]),
    .b(al_f2330f79[11]),
    .c(al_18077581[31]),
    .d(al_18077581[11]),
    .o(al_168e1cf3));
  AL_MAP_LUT6 #(
    .EQN("(B*A*(F@D)*(E@C))"),
    .INIT(64'h0008008008008000))
    al_c36dd5cd (
    .a(al_e2608c20),
    .b(al_168e1cf3),
    .c(al_f2330f79[27]),
    .d(al_f2330f79[15]),
    .e(al_18077581[27]),
    .f(al_18077581[15]),
    .o(al_2c27d715));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_a54e6d34 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[28]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_3b8c31d7),
    .o(al_f2330f79[28]));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    al_b1a5c121 (
    .a(al_f2330f79[18]),
    .b(al_f2330f79[9]),
    .c(al_18077581[18]),
    .d(al_18077581[9]),
    .o(al_6631dfe9));
  AL_MAP_LUT6 #(
    .EQN("(B*A*(F@D)*(E@C))"),
    .INIT(64'h0008008008008000))
    al_4cf6a0a3 (
    .a(al_2c27d715),
    .b(al_6631dfe9),
    .c(al_f2330f79[29]),
    .d(al_f2330f79[26]),
    .e(al_18077581[29]),
    .f(al_18077581[26]),
    .o(al_f3435a5b));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    al_3c91d255 (
    .a(al_f2330f79[19]),
    .b(al_f2330f79[5]),
    .c(al_18077581[19]),
    .d(al_18077581[5]),
    .o(al_cdd52893));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@C)*(D@B))"),
    .INIT(32'h02082080))
    al_f2d201d2 (
    .a(al_cdd52893),
    .b(al_f2330f79[17]),
    .c(al_f2330f79[12]),
    .d(al_18077581[17]),
    .e(al_18077581[12]),
    .o(al_626d1d9f));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@C)*(D@B))"),
    .INIT(32'h02082080))
    al_ecc85b60 (
    .a(al_626d1d9f),
    .b(al_f2330f79[21]),
    .c(al_f2330f79[10]),
    .d(al_18077581[21]),
    .e(al_18077581[10]),
    .o(al_ad3403a8));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_503a135d (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[27]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_102b7ad2),
    .o(al_f2330f79[27]));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    al_7912b7c2 (
    .a(al_f2330f79[8]),
    .b(al_f2330f79[7]),
    .c(al_18077581[7]),
    .d(al_18077581[8]),
    .o(al_faa08495));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@C)*(D@B))"),
    .INIT(32'h02082080))
    al_770fcb5d (
    .a(al_faa08495),
    .b(al_f2330f79[28]),
    .c(al_f2330f79[20]),
    .d(al_18077581[28]),
    .e(al_18077581[20]),
    .o(al_4580e6f4));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    al_6ded938d (
    .a(al_f2330f79[13]),
    .b(al_f2330f79[6]),
    .c(al_18077581[13]),
    .d(al_18077581[6]),
    .o(al_5b3bb87e));
  AL_MAP_LUT6 #(
    .EQN("(B*A*(F@D)*(E@C))"),
    .INIT(64'h0008008008008000))
    al_1c6ba0de (
    .a(al_4580e6f4),
    .b(al_5b3bb87e),
    .c(al_f2330f79[30]),
    .d(al_f2330f79[14]),
    .e(al_18077581[30]),
    .f(al_18077581[14]),
    .o(al_5c333c82));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    al_e8fb522a (
    .a(al_f2330f79[23]),
    .b(al_f2330f79[22]),
    .c(al_18077581[23]),
    .d(al_18077581[22]),
    .o(al_8e80a953));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_5ae3117a (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[26]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_6ec45564),
    .o(al_f2330f79[26]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@C)*(D@B))"),
    .INIT(32'h02082080))
    al_7cc6f9c3 (
    .a(al_8e80a953),
    .b(al_f2330f79[24]),
    .c(al_f2330f79[16]),
    .d(al_18077581[24]),
    .e(al_18077581[16]),
    .o(al_43f03d72));
  AL_MAP_LUT6 #(
    .EQN("((D@C)*(E@B)*(F@A))"),
    .INIT(64'h0110044002200880))
    al_60701873 (
    .a(al_f2330f79[4]),
    .b(al_f2330f79[2]),
    .c(al_f2330f79[1]),
    .d(al_18077581[1]),
    .e(al_18077581[2]),
    .f(al_18077581[4]),
    .o(al_13e18942));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_1fbba009 (
    .a(al_f3435a5b),
    .b(al_ad3403a8),
    .c(al_5c333c82),
    .d(al_43f03d72),
    .e(al_13e18942),
    .o(al_bdade024));
  AL_MAP_LUT6 #(
    .EQN("(D*(A*~(B)*~(C)*~(E)*~(F)+A*B*~(C)*~(E)*~(F)+~(A)*~(B)*C*~(E)*~(F)+~(A)*B*C*~(E)*~(F)+~(A)*B*~(C)*E*~(F)+A*B*~(C)*E*~(F)+~(A)*B*C*E*~(F)+A*B*C*E*~(F)+~(A)*B*~(C)*~(E)*F+A*B*~(C)*~(E)*F+~(A)*~(B)*C*~(E)*F+A*~(B)*C*~(E)*F+~(A)*B*~(C)*E*F+A*B*~(C)*E*F+~(A)*~(B)*C*E*F+A*~(B)*C*E*F))"),
    .INIT(64'h3c003c00cc005a00))
    al_862e1c4 (
    .a(al_bdade024),
    .b(al_eebab250),
    .c(al_bb6625de[1]),
    .d(al_580ff8b7[0]),
    .e(dBusAhb_HSIZE[1]),
    .f(al_e03b3126[14]),
    .o(al_b380555));
  AL_MAP_LUT3 #(
    .EQN("~(B@(~C*~A))"),
    .INIT(8'h36))
    al_8418a653 (
    .a(al_b380555),
    .b(al_86fb87b9),
    .c(al_580ff8b7[1]),
    .o(al_4357844d));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_d8c6789e (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[25]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_e611ec68),
    .o(al_f2330f79[25]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_fdb46626 (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[24]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_53b3dbc6),
    .o(al_f2330f79[24]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3550355f))
    al_d952893f (
    .a(al_e03b3126[31]),
    .b(al_9bf95cff[23]),
    .c(al_a1e88c0c[0]),
    .d(al_a1e88c0c[1]),
    .e(al_1f5093b5),
    .o(al_f2330f79[23]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ad9d68d5 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[0]),
    .d(al_1891b3c7),
    .o(al_d57349d9[0]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_71b0074d (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[10]),
    .d(al_407c8ac1),
    .o(al_d57349d9[10]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_dfcfd6f8 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[11]),
    .d(al_fdf9f0dc),
    .o(al_d57349d9[11]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_793c0a85 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[12]),
    .d(al_b5bf2603),
    .o(al_d57349d9[12]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_f2cca1bc (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[13]),
    .d(al_c8ba6c61),
    .o(al_d57349d9[13]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_51717195 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[14]),
    .d(al_59be2ab1),
    .o(al_d57349d9[14]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_70c2c38a (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[15]),
    .d(al_8488923),
    .o(al_d57349d9[15]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_c0fa6af6 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[16]),
    .d(al_5727b773),
    .o(al_d57349d9[16]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_db372661 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[17]),
    .d(al_eead7739),
    .o(al_d57349d9[17]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_c3956698 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[18]),
    .d(al_f430a5aa),
    .o(al_d57349d9[18]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_a470c15c (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[19]),
    .d(al_cd498e9f),
    .o(al_d57349d9[19]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_3a1802d6 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[1]),
    .d(al_512b1421),
    .o(al_d57349d9[1]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_1c5b45e7 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[20]),
    .d(al_3656d228),
    .o(al_d57349d9[20]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_59a0ec9b (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[21]),
    .d(al_30f08f9c),
    .o(al_d57349d9[21]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_43c9860b (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[22]),
    .d(al_bf6a3977),
    .o(al_d57349d9[22]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_c5b9b485 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[23]),
    .d(al_2ede456b),
    .o(al_d57349d9[23]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ec94f337 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[24]),
    .d(al_3a7c5a5),
    .o(al_d57349d9[24]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_4d40a601 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[25]),
    .d(al_9b707062),
    .o(al_d57349d9[25]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_80ac2233 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[26]),
    .d(al_a69cec28),
    .o(al_d57349d9[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ed3af229 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[27]),
    .d(al_d78f6bd4),
    .o(al_d57349d9[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_e309daac (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[28]),
    .d(al_cae21d2e),
    .o(al_d57349d9[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_56d9993f (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[29]),
    .d(al_19c0990d),
    .o(al_d57349d9[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_cb5b2781 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[2]),
    .d(al_80e2c141),
    .o(al_d57349d9[2]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_7b6dd4e9 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[30]),
    .d(al_cacb44c4),
    .o(al_d57349d9[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_74fa3473 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[31]),
    .d(al_14b732b9),
    .o(al_d57349d9[31]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_80c127a6 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[3]),
    .d(al_1e979a01),
    .o(al_d57349d9[3]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_b109d359 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[4]),
    .d(al_5df930ee),
    .o(al_d57349d9[4]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_fd3db5a1 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[5]),
    .d(al_8e267e24),
    .o(al_d57349d9[5]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_e2f532ce (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[6]),
    .d(al_e163f204),
    .o(al_d57349d9[6]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_9a431603 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[7]),
    .d(al_a6e0ed04),
    .o(al_d57349d9[7]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_b94f3f86 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[8]),
    .d(al_a35cf148),
    .o(al_d57349d9[8]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_49957be0 (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_9bf95cff[9]),
    .d(al_728c73ac),
    .o(al_d57349d9[9]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_8e999b1c (
    .a(al_580ff8b7[0]),
    .b(al_580ff8b7[1]),
    .c(al_e03b3126[20]),
    .o(al_35295e0a[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*B)))"),
    .INIT(16'hd500))
    al_4d95c81d (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[30]),
    .o(al_35295e0a[10]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hd5d0c5c015100500))
    al_d0b77bf0 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[7]),
    .e(al_e03b3126[20]),
    .f(al_e03b3126[31]),
    .o(al_35295e0a[11]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf4550400))
    al_f1d1937c (
    .a(al_86fb87b9),
    .b(al_bb6625de[1]),
    .c(al_580ff8b7[0]),
    .d(al_580ff8b7[1]),
    .e(al_e03b3126[31]),
    .o(al_35295e0a[12]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5c51000))
    al_4d8a37a4 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(dBusAhb_HSIZE[1]),
    .e(al_e03b3126[31]),
    .o(al_35295e0a[13]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5c51000))
    al_238cb3df (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[14]),
    .e(al_e03b3126[31]),
    .o(al_35295e0a[14]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5c51000))
    al_a277553f (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[15]),
    .e(al_e03b3126[31]),
    .o(al_35295e0a[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5c51000))
    al_b3c1ce97 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[16]),
    .e(al_e03b3126[31]),
    .o(al_35295e0a[16]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5c51000))
    al_865b8be6 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[17]),
    .e(al_e03b3126[31]),
    .o(al_35295e0a[17]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5c51000))
    al_f1326a29 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[18]),
    .e(al_e03b3126[31]),
    .o(al_35295e0a[18]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5c51000))
    al_81d0c639 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[19]),
    .e(al_e03b3126[31]),
    .o(al_35295e0a[19]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfbbbfb8808bb0888))
    al_b1fa0a44 (
    .a(al_9bcd349b),
    .b(al_86fb87b9),
    .c(al_580ff8b7[0]),
    .d(al_580ff8b7[1]),
    .e(al_e03b3126[8]),
    .f(al_e03b3126[21]),
    .o(al_35295e0a[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*B)))"),
    .INIT(16'hd500))
    al_40e30717 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[31]),
    .o(al_35295e0a[20]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf777f74404770444))
    al_b02eebe2 (
    .a(al_9bcd349b),
    .b(al_86fb87b9),
    .c(al_580ff8b7[0]),
    .d(al_580ff8b7[1]),
    .e(al_e03b3126[9]),
    .f(al_e03b3126[22]),
    .o(al_35295e0a[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5d00500))
    al_ddc7bada (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[10]),
    .e(al_e03b3126[23]),
    .o(al_35295e0a[3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hd5d00500))
    al_49d8fa44 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[11]),
    .e(al_e03b3126[24]),
    .o(al_35295e0a[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*B)))"),
    .INIT(16'hd500))
    al_6abecd22 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[25]),
    .o(al_35295e0a[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*B)))"),
    .INIT(16'hd500))
    al_27217297 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[26]),
    .o(al_35295e0a[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*B)))"),
    .INIT(16'hd500))
    al_dfa05d12 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[27]),
    .o(al_35295e0a[7]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*B)))"),
    .INIT(16'hd500))
    al_366ff128 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[28]),
    .o(al_35295e0a[8]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*B)))"),
    .INIT(16'hd500))
    al_5a968ec3 (
    .a(al_86fb87b9),
    .b(al_580ff8b7[0]),
    .c(al_580ff8b7[1]),
    .d(al_e03b3126[29]),
    .o(al_35295e0a[9]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*~C*B*~A)"),
    .INIT(64'h0400000000000000))
    al_780062b9 (
    .a(al_85a2bdb0[23]),
    .b(al_85a2bdb0[24]),
    .c(al_85a2bdb0[25]),
    .d(al_85a2bdb0[29]),
    .e(al_85a2bdb0[30]),
    .f(al_85a2bdb0[31]),
    .o(al_c36f1efd));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*~C*B*~A)"),
    .INIT(64'h0000000400000000))
    al_11a4a5e1 (
    .a(al_85a2bdb0[20]),
    .b(al_85a2bdb0[21]),
    .c(al_85a2bdb0[22]),
    .d(al_85a2bdb0[26]),
    .e(al_85a2bdb0[27]),
    .f(al_85a2bdb0[28]),
    .o(al_6f3fdf2e));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_14a7fd97 (
    .a(al_c36f1efd),
    .b(al_6f3fdf2e),
    .o(al_82a1cc96));
  AL_DFF_X al_3c443a3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_82a1cc96),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_235de557));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_7135b43f (
    .a(al_c281f5b2),
    .b(al_a4b1734c),
    .c(al_85a2bdb0[20]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[22]),
    .o(al_163b1f63));
  AL_DFF_X al_36516a94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_163b1f63),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e9897485));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_a1e13a9d (
    .a(al_c281f5b2),
    .b(al_a4b1734c),
    .c(al_85a2bdb0[20]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[22]),
    .o(al_dc7b4f80));
  AL_DFF_X al_b7ade031 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_dc7b4f80),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c55c5c3));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    al_90fd27e9 (
    .a(al_c281f5b2),
    .b(al_a4b1734c),
    .c(al_85a2bdb0[20]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[22]),
    .o(al_49e80206));
  AL_DFF_X al_17f23198 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_49e80206),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_804ebeec));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*~A)"),
    .INIT(64'h0000000000001000))
    al_922dde6a (
    .a(al_85a2bdb0[26]),
    .b(al_85a2bdb0[27]),
    .c(al_85a2bdb0[28]),
    .d(al_85a2bdb0[29]),
    .e(al_85a2bdb0[30]),
    .f(al_85a2bdb0[31]),
    .o(al_c281f5b2));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    al_a5a33452 (
    .a(al_c281f5b2),
    .b(al_a4b1734c),
    .c(al_85a2bdb0[20]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[22]),
    .o(al_4bc88254));
  AL_DFF_X al_f6a97a39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_4bc88254),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d19b9f6b));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_92b5fa6a (
    .a(al_d26be51c),
    .b(al_a4b1734c),
    .c(al_85a2bdb0[20]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[22]),
    .o(al_6782a2e8));
  AL_DFF_X al_7737ba74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6782a2e8),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8ea5e1));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    al_8da6f5f5 (
    .a(al_d26be51c),
    .b(al_a4b1734c),
    .c(al_85a2bdb0[20]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[22]),
    .o(al_58fb1503));
  AL_DFF_X al_a8258a6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_58fb1503),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4cc0b8dd));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_940b62ea (
    .a(al_85a2bdb0[23]),
    .b(al_85a2bdb0[24]),
    .c(al_85a2bdb0[25]),
    .o(al_a4b1734c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_2e08d759 (
    .a(al_85a2bdb0[26]),
    .b(al_85a2bdb0[27]),
    .c(al_85a2bdb0[28]),
    .d(al_85a2bdb0[29]),
    .e(al_85a2bdb0[30]),
    .f(al_85a2bdb0[31]),
    .o(al_d26be51c));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    al_c5a435af (
    .a(al_d26be51c),
    .b(al_a4b1734c),
    .c(al_85a2bdb0[20]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[22]),
    .o(al_895aceff));
  AL_DFF_X al_acb941a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_895aceff),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7610b7fc));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    al_9281d647 (
    .a(al_d26be51c),
    .b(al_a4b1734c),
    .c(al_85a2bdb0[20]),
    .d(al_85a2bdb0[21]),
    .e(al_85a2bdb0[22]),
    .o(al_709aaff2));
  AL_DFF_X al_f0ce852f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_709aaff2),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_809b319));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    al_c7a664f5 (
    .a(al_4d82afcf),
    .b(al_6893b11d),
    .o(al_cf7a2555));
  AL_DFF_X al_22265819 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf7a2555),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bb6ca07d));
  AL_MAP_LUT3 #(
    .EQN("(C*(B@A))"),
    .INIT(8'h60))
    al_ecbbf12e (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_14b732b9),
    .o(al_da34572b[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_a0a0c442 (
    .a(al_bb6625de[1]),
    .b(dBusAhb_HSIZE[1]),
    .c(al_60dd36d7),
    .o(al_65e3dd93[16]));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8f3029b1 (
    .i(al_8074bdb[0]),
    .o(al_3e08733b[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e81abc87 (
    .i(al_3e08733b[0]),
    .o(al_1891b3c7));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_955407d4 (
    .i(al_8074bdb[10]),
    .o(al_3e08733b[10]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_8af3d71d (
    .i(al_3e08733b[10]),
    .o(al_407c8ac1));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c9c7d14b (
    .i(al_8074bdb[11]),
    .o(al_3e08733b[11]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_120af05b (
    .i(al_3e08733b[11]),
    .o(al_fdf9f0dc));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_19720074 (
    .i(al_8074bdb[12]),
    .o(al_3e08733b[12]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_8c001ff7 (
    .i(al_3e08733b[12]),
    .o(al_b5bf2603));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5fc0cd55 (
    .i(al_8074bdb[13]),
    .o(al_3e08733b[13]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_37d9b9ce (
    .i(al_3e08733b[13]),
    .o(al_c8ba6c61));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b01d91c4 (
    .i(al_8074bdb[14]),
    .o(al_3e08733b[14]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c8abb69c (
    .i(al_3e08733b[14]),
    .o(al_59be2ab1));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_caa54e6a (
    .i(al_8074bdb[15]),
    .o(al_3e08733b[15]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_340580 (
    .i(al_3e08733b[15]),
    .o(al_8488923));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4b9b2c41 (
    .i(al_8074bdb[16]),
    .o(al_3e08733b[16]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9449a325 (
    .i(al_3e08733b[16]),
    .o(al_5727b773));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7cbe8a33 (
    .i(al_8074bdb[17]),
    .o(al_3e08733b[17]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_14ae075f (
    .i(al_3e08733b[17]),
    .o(al_eead7739));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_dd686d2a (
    .i(al_8074bdb[18]),
    .o(al_3e08733b[18]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_36c6aea1 (
    .i(al_3e08733b[18]),
    .o(al_f430a5aa));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_adb56be5 (
    .i(al_8074bdb[19]),
    .o(al_3e08733b[19]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c1ddb63d (
    .i(al_3e08733b[19]),
    .o(al_cd498e9f));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_aafbf6e4 (
    .i(al_8074bdb[1]),
    .o(al_3e08733b[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_28037775 (
    .i(al_3e08733b[1]),
    .o(al_512b1421));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_7fa7f638 (
    .i(al_8074bdb[20]),
    .o(al_3e08733b[20]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3d96e342 (
    .i(al_3e08733b[20]),
    .o(al_3656d228));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1a327526 (
    .i(al_8074bdb[21]),
    .o(al_3e08733b[21]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9fd5fed0 (
    .i(al_3e08733b[21]),
    .o(al_30f08f9c));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_454f924e (
    .i(al_8074bdb[22]),
    .o(al_3e08733b[22]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_93f6269b (
    .i(al_3e08733b[22]),
    .o(al_bf6a3977));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_81d4ccad (
    .i(al_8074bdb[23]),
    .o(al_3e08733b[23]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_fecbe189 (
    .i(al_3e08733b[23]),
    .o(al_2ede456b));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8e64a90e (
    .i(al_8074bdb[24]),
    .o(al_3e08733b[24]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a1193750 (
    .i(al_3e08733b[24]),
    .o(al_3a7c5a5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_db1f6c12 (
    .i(al_8074bdb[25]),
    .o(al_3e08733b[25]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_3c598ccf (
    .i(al_3e08733b[25]),
    .o(al_9b707062));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d9b33f67 (
    .i(al_8074bdb[26]),
    .o(al_3e08733b[26]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_ab1bc58e (
    .i(al_3e08733b[26]),
    .o(al_a69cec28));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3cf24ecc (
    .i(al_8074bdb[27]),
    .o(al_3e08733b[27]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d41eae05 (
    .i(al_3e08733b[27]),
    .o(al_d78f6bd4));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f3ec7d81 (
    .i(al_8074bdb[28]),
    .o(al_3e08733b[28]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d2630ace (
    .i(al_3e08733b[28]),
    .o(al_cae21d2e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_59f3e7fd (
    .i(al_8074bdb[29]),
    .o(al_3e08733b[29]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_7183c019 (
    .i(al_3e08733b[29]),
    .o(al_19c0990d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_17f9e732 (
    .i(al_8074bdb[2]),
    .o(al_3e08733b[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b9cbbaf6 (
    .i(al_3e08733b[2]),
    .o(al_80e2c141));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f4b686d9 (
    .i(al_8074bdb[30]),
    .o(al_3e08733b[30]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_48497b90 (
    .i(al_3e08733b[30]),
    .o(al_cacb44c4));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_dd533a9b (
    .i(al_8074bdb[31]),
    .o(al_3e08733b[31]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_722f41f8 (
    .i(al_3e08733b[31]),
    .o(al_14b732b9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_577e6634 (
    .i(al_8074bdb[3]),
    .o(al_3e08733b[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_75e97d68 (
    .i(al_3e08733b[3]),
    .o(al_1e979a01));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_bfe0ce41 (
    .i(al_8074bdb[4]),
    .o(al_3e08733b[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_75e08010 (
    .i(al_3e08733b[4]),
    .o(al_5df930ee));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_6ff4544c (
    .i(al_8074bdb[5]),
    .o(al_3e08733b[5]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_c023be93 (
    .i(al_3e08733b[5]),
    .o(al_8e267e24));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_67a0c20f (
    .i(al_8074bdb[6]),
    .o(al_3e08733b[6]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9eb63343 (
    .i(al_3e08733b[6]),
    .o(al_e163f204));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_18337bbe (
    .i(al_8074bdb[7]),
    .o(al_3e08733b[7]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e3d06bd9 (
    .i(al_3e08733b[7]),
    .o(al_a6e0ed04));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4caea158 (
    .i(al_8074bdb[8]),
    .o(al_3e08733b[8]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e262f530 (
    .i(al_3e08733b[8]),
    .o(al_a35cf148));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_54ccdb82 (
    .i(al_8074bdb[9]),
    .o(al_3e08733b[9]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b1c1d3b9 (
    .i(al_3e08733b[9]),
    .o(al_728c73ac));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8c38761f (
    .i(al_2f7928e2[0]),
    .o(al_b541ca02[0]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4981840d (
    .i(al_b541ca02[0]),
    .o(al_f4b5275b));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_a72f763a (
    .i(al_2f7928e2[10]),
    .o(al_b541ca02[10]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_8ff0982c (
    .i(al_b541ca02[10]),
    .o(al_98804c07));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_78769376 (
    .i(al_2f7928e2[11]),
    .o(al_b541ca02[11]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_cfd5ee74 (
    .i(al_b541ca02[11]),
    .o(al_3ebb68c3));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_90e341a (
    .i(al_2f7928e2[12]),
    .o(al_b541ca02[12]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d1af3d15 (
    .i(al_b541ca02[12]),
    .o(al_d00a6f56));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8266c23c (
    .i(al_2f7928e2[13]),
    .o(al_b541ca02[13]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6123a27c (
    .i(al_b541ca02[13]),
    .o(al_e6455839));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f8959082 (
    .i(al_2f7928e2[14]),
    .o(al_b541ca02[14]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_620376c (
    .i(al_b541ca02[14]),
    .o(al_7e6320f4));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_8d3cbc3c (
    .i(al_2f7928e2[15]),
    .o(al_b541ca02[15]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_dba4b264 (
    .i(al_b541ca02[15]),
    .o(al_f61ec828));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_66e382fb (
    .i(al_2f7928e2[16]),
    .o(al_b541ca02[16]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6bbed6e9 (
    .i(al_b541ca02[16]),
    .o(al_7d27d680));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_871fa1c0 (
    .i(al_2f7928e2[17]),
    .o(al_b541ca02[17]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_f5fda335 (
    .i(al_b541ca02[17]),
    .o(al_d76255c5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_521f14f0 (
    .i(al_2f7928e2[18]),
    .o(al_b541ca02[18]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_475b879d (
    .i(al_b541ca02[18]),
    .o(al_3b0f4da7));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_cddd8744 (
    .i(al_2f7928e2[19]),
    .o(al_b541ca02[19]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_fe64d223 (
    .i(al_b541ca02[19]),
    .o(al_c7df4b4d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_3e85601f (
    .i(al_2f7928e2[1]),
    .o(al_b541ca02[1]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b10558cf (
    .i(al_b541ca02[1]),
    .o(al_2370214));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d8f89c16 (
    .i(al_2f7928e2[20]),
    .o(al_b541ca02[20]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d60ea349 (
    .i(al_b541ca02[20]),
    .o(al_a831c176));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_16733456 (
    .i(al_2f7928e2[21]),
    .o(al_b541ca02[21]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_322a1e3e (
    .i(al_b541ca02[21]),
    .o(al_658bb789));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_88acddee (
    .i(al_2f7928e2[22]),
    .o(al_b541ca02[22]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_d00a514a (
    .i(al_b541ca02[22]),
    .o(al_ffc4fe26));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1fdead20 (
    .i(al_2f7928e2[23]),
    .o(al_b541ca02[23]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_65ef3db2 (
    .i(al_b541ca02[23]),
    .o(al_1f5093b5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_c886e514 (
    .i(al_2f7928e2[24]),
    .o(al_b541ca02[24]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b87e3e22 (
    .i(al_b541ca02[24]),
    .o(al_53b3dbc6));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_4a4a7846 (
    .i(al_2f7928e2[25]),
    .o(al_b541ca02[25]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_9dc296e5 (
    .i(al_b541ca02[25]),
    .o(al_e611ec68));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_f37418b0 (
    .i(al_2f7928e2[26]),
    .o(al_b541ca02[26]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_4b8db41d (
    .i(al_b541ca02[26]),
    .o(al_6ec45564));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_86347ae (
    .i(al_2f7928e2[27]),
    .o(al_b541ca02[27]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_2af0c0cc (
    .i(al_b541ca02[27]),
    .o(al_102b7ad2));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_5ff7c132 (
    .i(al_2f7928e2[28]),
    .o(al_b541ca02[28]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_a1e1f3cb (
    .i(al_b541ca02[28]),
    .o(al_3b8c31d7));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1f80388f (
    .i(al_2f7928e2[29]),
    .o(al_b541ca02[29]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_aabc6c2c (
    .i(al_b541ca02[29]),
    .o(al_3626cb0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ea537ff (
    .i(al_2f7928e2[2]),
    .o(al_b541ca02[2]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_ef55ecd (
    .i(al_b541ca02[2]),
    .o(al_bf952132));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_bf437fcb (
    .i(al_2f7928e2[30]),
    .o(al_b541ca02[30]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_f2183da5 (
    .i(al_b541ca02[30]),
    .o(al_f1bb92e9));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_b44f4bb4 (
    .i(al_2f7928e2[31]),
    .o(al_b541ca02[31]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_ecccbf64 (
    .i(al_b541ca02[31]),
    .o(al_60dd36d7));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_ad861c1f (
    .i(al_2f7928e2[3]),
    .o(al_b541ca02[3]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_e963a1b7 (
    .i(al_b541ca02[3]),
    .o(al_76a52f3d));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_768e2602 (
    .i(al_2f7928e2[4]),
    .o(al_b541ca02[4]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_1759dc0e (
    .i(al_b541ca02[4]),
    .o(al_c861c8f0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_55942bd0 (
    .i(al_2f7928e2[5]),
    .o(al_b541ca02[5]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_791b8e1d (
    .i(al_b541ca02[5]),
    .o(al_8a841cb4));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_214bbafb (
    .i(al_2f7928e2[6]),
    .o(al_b541ca02[6]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_848a4298 (
    .i(al_b541ca02[6]),
    .o(al_33a2911e));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_1813be6a (
    .i(al_2f7928e2[7]),
    .o(al_b541ca02[7]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_b6f391ca (
    .i(al_b541ca02[7]),
    .o(al_73fb1ee5));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_d1813a77 (
    .i(al_2f7928e2[8]),
    .o(al_b541ca02[8]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_efc97415 (
    .i(al_b541ca02[8]),
    .o(al_bdb28b76));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    al_df34a017 (
    .i(al_2f7928e2[9]),
    .o(al_b541ca02[9]));
  AL_BUFKEEP #(
    .KEEP("IN"))
    al_6b6f3280 (
    .i(al_b541ca02[9]),
    .o(al_6d92b3c6));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    al_3974232d (
    .a(al_6a0e908c),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_e379ebb5),
    .o(al_592c9a6));
  AL_MAP_LUT6 #(
    .EQN("((F*B)*~((~E*D*A))*~(C)+(F*B)*(~E*D*A)*~(C)+~((F*B))*(~E*D*A)*C+(F*B)*(~E*D*A)*C)"),
    .INIT(64'h0c0cac0c0000a000))
    al_75eabd89 (
    .a(al_3f1d46e5),
    .b(al_592c9a6),
    .c(al_5a744f0f),
    .d(al_6f08d701),
    .e(al_f6cd735f),
    .f(al_523cde28),
    .o(al_7c88a272));
  AL_DFF_X al_78db16a (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_7c88a272),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_523cde28));
  AL_DFF_X al_10fe5e3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_7bc36116),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_673a4598));
  AL_DFF_X al_a9e0a4d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_4357844d),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd3d5e6f));
  AL_DFF_X al_47fce0dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6b2d5c80),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cdace779));
  AL_DFF_X al_a97757a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c5b8f9ea),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b2739b77));
  AL_DFF_X al_c839841e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9a05e7eb),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3290619));
  AL_DFF_X al_4bcd89cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32fedef4),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e3edcf1a));
  AL_DFF_X al_ac8b4578 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HWRITE),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_587b9831));
  AL_DFF_X al_db3d0849 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_44595135),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24641d37));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_b2f3fb9 (
    .a(al_e108f0ff[0]),
    .b(al_e108f0ff[3]),
    .c(al_e108f0ff[5]),
    .d(al_d264c8ee[0]),
    .e(al_d264c8ee[3]),
    .f(al_d264c8ee[5]),
    .o(al_691a2d0a));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(E*B)*~(D*A))"),
    .INIT(64'h0103050f113355ff))
    al_431ebf6b (
    .a(al_e108f0ff[1]),
    .b(al_e108f0ff[2]),
    .c(al_e108f0ff[4]),
    .d(al_d264c8ee[1]),
    .e(al_d264c8ee[2]),
    .f(al_d264c8ee[4]),
    .o(al_4f8cc1b7));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    al_d590b9e5 (
    .a(al_691a2d0a),
    .b(al_4f8cc1b7),
    .o(al_abe3d564));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_1fe38e43 (
    .a(al_a3de3eda[0]),
    .b(al_a3de3eda[1]),
    .c(al_a3de3eda[2]),
    .d(al_a3de3eda[3]),
    .o(al_a44ada9e));
  AL_DFF_X al_74473634 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(CORE_TDI),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2802ceac));
  AL_DFF_X al_d3c490c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_56c9e07a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5356e8f));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf753229d))
    al_9f24e20e (
    .a(CORE_TMS),
    .b(al_549b2fd9[0]),
    .c(al_549b2fd9[1]),
    .d(al_549b2fd9[2]),
    .e(al_549b2fd9[3]),
    .o(al_53f57cc3[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h3a5c3410))
    al_42b6b64e (
    .a(CORE_TMS),
    .b(al_549b2fd9[0]),
    .c(al_549b2fd9[1]),
    .d(al_549b2fd9[2]),
    .e(al_549b2fd9[3]),
    .o(al_53f57cc3[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h2fa077c0))
    al_7641fe4b (
    .a(CORE_TMS),
    .b(al_549b2fd9[0]),
    .c(al_549b2fd9[1]),
    .d(al_549b2fd9[2]),
    .e(al_549b2fd9[3]),
    .o(al_53f57cc3[2]));
  AL_MAP_LUT5 #(
    .EQN("(A*B*~(C)*~(D)*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hbff68808))
    al_40e1f2a7 (
    .a(CORE_TMS),
    .b(al_549b2fd9[0]),
    .c(al_549b2fd9[1]),
    .d(al_549b2fd9[2]),
    .e(al_549b2fd9[3]),
    .o(al_53f57cc3[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_30b9de28 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[0]),
    .d(al_d48366e1[1]),
    .e(al_a45b58d1),
    .o(al_8eb7c3ef[0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_97bfa6f7 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[10]),
    .d(al_d48366e1[11]),
    .e(al_156dfeae[8]),
    .o(al_8eb7c3ef[10]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_3f25f308 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[11]),
    .d(al_d48366e1[12]),
    .e(al_156dfeae[9]),
    .o(al_8eb7c3ef[11]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_ad047a7b (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[12]),
    .d(al_d48366e1[13]),
    .e(al_156dfeae[10]),
    .o(al_8eb7c3ef[12]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_9e9ac1a6 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[13]),
    .d(al_d48366e1[14]),
    .e(al_156dfeae[11]),
    .o(al_8eb7c3ef[13]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_292064a1 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[14]),
    .d(al_d48366e1[15]),
    .e(al_156dfeae[12]),
    .o(al_8eb7c3ef[14]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_437a2474 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[15]),
    .d(al_d48366e1[16]),
    .e(al_156dfeae[13]),
    .o(al_8eb7c3ef[15]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_5a5c3ba1 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[16]),
    .d(al_d48366e1[17]),
    .e(al_156dfeae[14]),
    .o(al_8eb7c3ef[16]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_adebddc6 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[17]),
    .d(al_d48366e1[18]),
    .e(al_156dfeae[15]),
    .o(al_8eb7c3ef[17]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_b56da512 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[18]),
    .d(al_d48366e1[19]),
    .e(al_156dfeae[16]),
    .o(al_8eb7c3ef[18]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_cb1e6f3 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[19]),
    .d(al_d48366e1[20]),
    .e(al_156dfeae[17]),
    .o(al_8eb7c3ef[19]));
  AL_MAP_LUT4 #(
    .EQN("((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'hdc10))
    al_f363e6fc (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[1]),
    .d(al_d48366e1[2]),
    .o(al_8eb7c3ef[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_a7d19917 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[20]),
    .d(al_d48366e1[21]),
    .e(al_156dfeae[18]),
    .o(al_8eb7c3ef[20]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_cc7447d8 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[21]),
    .d(al_d48366e1[22]),
    .e(al_156dfeae[19]),
    .o(al_8eb7c3ef[21]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_f8e42e00 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[22]),
    .d(al_d48366e1[23]),
    .e(al_156dfeae[20]),
    .o(al_8eb7c3ef[22]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_b6ac5ba9 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[23]),
    .d(al_d48366e1[24]),
    .e(al_156dfeae[21]),
    .o(al_8eb7c3ef[23]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_7b236ff4 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[24]),
    .d(al_d48366e1[25]),
    .e(al_156dfeae[22]),
    .o(al_8eb7c3ef[24]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_dcda6aa0 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[25]),
    .d(al_d48366e1[26]),
    .e(al_156dfeae[23]),
    .o(al_8eb7c3ef[25]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_818971b1 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[26]),
    .d(al_d48366e1[27]),
    .e(al_156dfeae[24]),
    .o(al_8eb7c3ef[26]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_1214521c (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[27]),
    .d(al_d48366e1[28]),
    .e(al_156dfeae[25]),
    .o(al_8eb7c3ef[27]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_adaa600c (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[28]),
    .d(al_d48366e1[29]),
    .e(al_156dfeae[26]),
    .o(al_8eb7c3ef[28]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_387cf9e3 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[29]),
    .d(al_d48366e1[30]),
    .e(al_156dfeae[27]),
    .o(al_8eb7c3ef[29]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_7fc75ff1 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[2]),
    .d(al_d48366e1[3]),
    .e(al_156dfeae[0]),
    .o(al_8eb7c3ef[2]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_d219fe8c (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[30]),
    .d(al_d48366e1[31]),
    .e(al_156dfeae[28]),
    .o(al_8eb7c3ef[30]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    al_d34f3f5c (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .o(al_a4860493));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_345afd13 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[31]),
    .d(al_d48366e1[32]),
    .e(al_156dfeae[29]),
    .o(al_8eb7c3ef[31]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_a46b9e77 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[32]),
    .d(al_d48366e1[33]),
    .e(al_156dfeae[30]),
    .o(al_8eb7c3ef[32]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_e583562c (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(CORE_TDI),
    .d(al_d48366e1[33]),
    .e(al_156dfeae[31]),
    .o(al_8eb7c3ef[33]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_e13e8779 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[3]),
    .d(al_d48366e1[4]),
    .e(al_156dfeae[1]),
    .o(al_8eb7c3ef[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_e15ebaad (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[4]),
    .d(al_d48366e1[5]),
    .e(al_156dfeae[2]),
    .o(al_8eb7c3ef[4]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_2d5bbc11 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[5]),
    .d(al_d48366e1[6]),
    .e(al_156dfeae[3]),
    .o(al_8eb7c3ef[5]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_eec15779 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[6]),
    .d(al_d48366e1[7]),
    .e(al_156dfeae[4]),
    .o(al_8eb7c3ef[6]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_99abec71 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[7]),
    .d(al_d48366e1[8]),
    .e(al_156dfeae[5]),
    .o(al_8eb7c3ef[7]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_4de26e5 (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[8]),
    .d(al_d48366e1[9]),
    .e(al_156dfeae[6]),
    .o(al_8eb7c3ef[8]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_f6c1078b (
    .a(al_a4860493),
    .b(al_f5a4c6e6),
    .c(al_d48366e1[9]),
    .d(al_d48366e1[10]),
    .e(al_156dfeae[7]),
    .o(al_8eb7c3ef[9]));
  AL_DFF_X al_f471f8d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8bf04ef0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_871b264a));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_717afbd3 (
    .a(al_2802ceac),
    .b(al_b5356e8f),
    .c(al_871b264a),
    .o(al_8bf04ef0));
  AL_DFF_X al_9490ddd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_b7e97af1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d7a8be80));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    al_3411eaca (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .o(al_f5a4c6e6));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_863ffdcc (
    .a(al_f5a4c6e6),
    .b(al_a3de3eda[0]),
    .c(al_a3de3eda[1]),
    .d(al_a3de3eda[2]),
    .e(al_a3de3eda[3]),
    .o(al_56c9e07a));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ede57c5 (
    .a(al_56c9e07a),
    .b(al_b5356e8f),
    .c(al_d7a8be80),
    .o(al_b7e97af1));
  AL_DFF_X al_3e99ad6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_13a562ab),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d28932f));
  AL_DFF_X al_3838b0a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6d28932f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eeed7a72));
  AL_DFF_0 al_b25d2722 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_4c35eef2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13a562ab));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e5716b76 (
    .a(al_b5356e8f),
    .b(al_13a562ab),
    .o(al_4c35eef2));
  AL_DFF_X al_b614f99c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_59c9e271),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2ae0151));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b5bbabfe (
    .a(al_c4f8cd6c),
    .b(al_871b264a),
    .c(al_c2ae0151),
    .o(al_59c9e271));
  AL_DFF_X al_d1e5efcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_31e2d17a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6380dbe7));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_8649d8d1 (
    .a(al_53ca6362),
    .b(al_eeed7a72),
    .o(al_c4f8cd6c));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b30e0cd9 (
    .a(al_c4f8cd6c),
    .b(al_d7a8be80),
    .c(al_6380dbe7),
    .o(al_31e2d17a));
  AL_DFF_X al_cdf4fd09 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c4f8cd6c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7b5abb5));
  AL_DFF_X al_efa9bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_eeed7a72),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53ca6362));
  AL_DFF_X al_95148300 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~CORE_TCK),
    .d(al_fa675d9c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(CORE_TDO));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_18d5aeae (
    .a(al_f5a4c6e6),
    .b(al_a3de3eda[0]),
    .c(al_a3de3eda[1]),
    .d(al_a3de3eda[2]),
    .e(al_a3de3eda[3]),
    .o(al_5c1a51fa));
  AL_DFF_X al_1c857cb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[8]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[8]));
  AL_DFF_X al_b6a60ff3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[9]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[9]));
  AL_DFF_X al_ed594fd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[10]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[10]));
  AL_DFF_X al_5bcb14ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[11]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[11]));
  AL_DFF_X al_6d78ff05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[12]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[12]));
  AL_DFF_X al_4a3c1d60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[13]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[13]));
  AL_DFF_X al_2bb5b87f (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[14]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[14]));
  AL_DFF_X al_4e091958 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[15]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[15]));
  AL_DFF_X al_88da4f8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[16]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[16]));
  AL_DFF_X al_5d24ee0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[17]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[17]));
  AL_DFF_X al_f603c107 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[0]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[0]));
  AL_DFF_X al_5c9a182 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[18]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[18]));
  AL_DFF_X al_a3e2566a (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[19]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[19]));
  AL_DFF_X al_d3b31986 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[20]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[20]));
  AL_DFF_X al_a7295b80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[21]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[21]));
  AL_DFF_X al_a6b380de (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[22]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[22]));
  AL_DFF_X al_72db48df (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[23]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[23]));
  AL_DFF_X al_50050383 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[24]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[24]));
  AL_DFF_X al_d1a4747 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[25]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[25]));
  AL_DFF_X al_654d6d9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[26]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[26]));
  AL_DFF_X al_6074b532 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[27]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[27]));
  AL_DFF_X al_659b2a2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[1]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[1]));
  AL_DFF_X al_5ec81828 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[28]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[28]));
  AL_DFF_X al_7ec51c7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[29]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[29]));
  AL_DFF_X al_39117b04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[30]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[30]));
  AL_DFF_X al_6dedc243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[31]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[31]));
  AL_DFF_X al_d9fa4ff8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[32]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[32]));
  AL_DFF_X al_7d4bfe86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[33]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[33]));
  AL_DFF_X al_c0328df5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[2]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[2]));
  AL_DFF_X al_a12aa5fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[3]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[3]));
  AL_DFF_X al_48f9b8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[4]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[4]));
  AL_DFF_X al_b1a59b72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[5]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[5]));
  AL_DFF_X al_269f950c (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[6]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[6]));
  AL_DFF_X al_4d4b88dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_8eb7c3ef[7]),
    .en(al_a44ada9e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d48366e1[7]));
  AL_DFF_X al_8a885193 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[9]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[8]));
  AL_DFF_X al_d4bf26a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[10]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[9]));
  AL_DFF_X al_aaa1dc97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[11]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[10]));
  AL_DFF_X al_f01dd73e (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[12]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[11]));
  AL_DFF_X al_74e99570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[13]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[12]));
  AL_DFF_X al_106721e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[14]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[13]));
  AL_DFF_X al_9ae735e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[15]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[14]));
  AL_DFF_X al_43f82305 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[16]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[15]));
  AL_DFF_X al_b577e5b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[17]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[16]));
  AL_DFF_X al_bd1d1fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[18]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[17]));
  AL_DFF_X al_a31d3527 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[1]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[0]));
  AL_DFF_X al_d1b26649 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[19]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[18]));
  AL_DFF_X al_3b79ab60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[20]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[19]));
  AL_DFF_X al_16e42d94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[21]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[20]));
  AL_DFF_X al_a0b67da9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[22]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[21]));
  AL_DFF_X al_11024e80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[23]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[22]));
  AL_DFF_X al_c24ca1b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[24]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[23]));
  AL_DFF_X al_d061eacf (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[25]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[24]));
  AL_DFF_X al_cbc78b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[26]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[25]));
  AL_DFF_X al_78fce76f (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[27]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[26]));
  AL_DFF_X al_d93f6ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[28]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[27]));
  AL_DFF_X al_cb487964 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[2]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[1]));
  AL_DFF_X al_de5e24d (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[29]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[28]));
  AL_DFF_X al_62709cab (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[30]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[29]));
  AL_DFF_X al_15e17adb (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[31]),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[30]));
  AL_DFF_X al_f4023da1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(CORE_TDI),
    .en(al_5c1a51fa),
    .sr(al_a4860493),
    .ss(1'b0),
    .q(al_a550c05f[31]));
  AL_DFF_X al_245e99b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[3]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[2]));
  AL_DFF_X al_41e2d963 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[4]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[3]));
  AL_DFF_X al_d60a83e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[5]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[4]));
  AL_DFF_X al_1b89e1c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[6]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[5]));
  AL_DFF_X al_3efe7213 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[7]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[6]));
  AL_DFF_X al_17bd2efd (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_a550c05f[8]),
    .en(al_5c1a51fa),
    .sr(1'b0),
    .ss(al_a4860493),
    .q(al_a550c05f[7]));
  AL_DFF_0 al_f0beebbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_53f57cc3[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_549b2fd9[0]));
  AL_DFF_0 al_880f05a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_53f57cc3[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_549b2fd9[1]));
  AL_DFF_0 al_2a248138 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_53f57cc3[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_549b2fd9[2]));
  AL_DFF_0 al_e22ce433 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_53f57cc3[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_549b2fd9[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*D*~(E)*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffbffe3f00800200))
    al_22d7a831 (
    .a(CORE_TDI),
    .b(al_549b2fd9[0]),
    .c(al_549b2fd9[1]),
    .d(al_549b2fd9[2]),
    .e(al_549b2fd9[3]),
    .f(al_a6bbd516[3]),
    .o(al_d9ff9b46));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffff0818f7ef0008))
    al_2f73eafd (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .e(al_a6bbd516[0]),
    .f(al_a6bbd516[1]),
    .o(al_ab1643c6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff70810f7e70000))
    al_d8e0a2fd (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .e(al_a6bbd516[1]),
    .f(al_a6bbd516[2]),
    .o(al_bc4322fc));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff70810f7e70000))
    al_f9222dbf (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .e(al_a6bbd516[2]),
    .f(al_a6bbd516[3]),
    .o(al_c3666229));
  AL_DFF_X al_b564218a (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_ab1643c6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6bbd516[0]));
  AL_DFF_X al_1d3bd47f (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_bc4322fc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6bbd516[1]));
  AL_DFF_X al_324d92cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_c3666229),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6bbd516[2]));
  AL_DFF_X al_bc879c15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_d9ff9b46),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6bbd516[3]));
  AL_DFF_X al_ec74a203 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_d72457d3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3de3eda[0]));
  AL_MAP_LUT6 #(
    .EQN("(F*~((E*D))*~((~C*~B*~A))+F*(E*D)*~((~C*~B*~A))+~(F)*(E*D)*(~C*~B*~A)+F*(E*D)*(~C*~B*~A))"),
    .INIT(64'hfffefefe01000000))
    al_7c560de2 (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .e(al_a6bbd516[3]),
    .f(al_a3de3eda[3]),
    .o(al_3d575f81));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~((~E*D))*~((~C*~B*~A))+~F*(~E*D)*~((~C*~B*~A))+~(~F)*(~E*D)*(~C*~B*~A)+~F*(~E*D)*(~C*~B*~A))"),
    .INIT(64'hfffffeff01010001))
    al_2daa9fb1 (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .e(al_a6bbd516[0]),
    .f(al_a3de3eda[0]),
    .o(al_d72457d3));
  AL_MAP_LUT6 #(
    .EQN("(F*~((E*D))*~((~C*~B*~A))+F*(E*D)*~((~C*~B*~A))+~(F)*(E*D)*(~C*~B*~A)+F*(E*D)*(~C*~B*~A))"),
    .INIT(64'hfffefefe01000000))
    al_e1125700 (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .e(al_a6bbd516[1]),
    .f(al_a3de3eda[1]),
    .o(al_9061aac4));
  AL_MAP_LUT6 #(
    .EQN("(F*~((E*D))*~((~C*~B*~A))+F*(E*D)*~((~C*~B*~A))+~(F)*(E*D)*(~C*~B*~A)+F*(E*D)*(~C*~B*~A))"),
    .INIT(64'hfffefefe01000000))
    al_de7bd908 (
    .a(al_549b2fd9[0]),
    .b(al_549b2fd9[1]),
    .c(al_549b2fd9[2]),
    .d(al_549b2fd9[3]),
    .e(al_a6bbd516[2]),
    .f(al_a3de3eda[2]),
    .o(al_ac066a39));
  AL_DFF_X al_89100783 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_9061aac4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3de3eda[1]));
  AL_DFF_X al_1d5792b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_ac066a39),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3de3eda[2]));
  AL_DFF_X al_81a1bb10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(CORE_TCK),
    .d(al_3d575f81),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3de3eda[3]));
  AL_DFF_X al_fe120d14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[8]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[8]));
  AL_DFF_X al_aa3c24f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[9]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[9]));
  AL_DFF_X al_e5fc30cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[10]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[10]));
  AL_DFF_X al_61f385e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[11]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[11]));
  AL_DFF_X al_c4fe8dfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[12]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[12]));
  AL_DFF_X al_a7521e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[13]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[13]));
  AL_DFF_X al_66547d20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[14]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[14]));
  AL_DFF_X al_7e48a106 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[15]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[15]));
  AL_DFF_X al_ae183d9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[16]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[16]));
  AL_DFF_X al_808e1a50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[17]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[17]));
  AL_DFF_X al_8ad3881e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_daece8d7[0]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[0]));
  AL_DFF_X al_710fedc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[18]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[18]));
  AL_DFF_X al_f55cf05b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[19]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[19]));
  AL_DFF_X al_f542ca28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[20]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[20]));
  AL_DFF_X al_a55cbc7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[21]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[21]));
  AL_DFF_X al_d6ec655d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[22]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[22]));
  AL_DFF_X al_3ada1a69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[23]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[23]));
  AL_DFF_X al_ddc0523e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[24]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[24]));
  AL_DFF_X al_4b4319f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[25]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[25]));
  AL_DFF_X al_23195ac7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[26]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[26]));
  AL_DFF_X al_e846f781 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[27]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[27]));
  AL_DFF_X al_2abc224b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_daece8d7[1]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[1]));
  AL_DFF_X al_612bfa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[28]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[28]));
  AL_DFF_X al_5a1c2a90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[29]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[29]));
  AL_DFF_X al_20ef96c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[30]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[30]));
  AL_DFF_X al_8c75e2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[31]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[31]));
  AL_DFF_X al_c4a7a267 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_daece8d7[2]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[2]));
  AL_DFF_X al_458abd37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_daece8d7[3]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[3]));
  AL_DFF_X al_391f9824 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_daece8d7[4]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[4]));
  AL_DFF_X al_8aac0a49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[5]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[5]));
  AL_DFF_X al_ab19853a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[6]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[6]));
  AL_DFF_X al_896cee58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_43722bf9[7]),
    .en(al_18c565c8),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_156dfeae[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_aa80ade7 (
    .a(al_d48366e1[0]),
    .b(al_a550c05f[0]),
    .c(al_a3de3eda[1]),
    .o(al_ee5ae3ff));
  AL_MAP_LUT6 #(
    .EQN("~(C*~((~F*~E*D*B))*~(A)+C*(~F*~E*D*B)*~(A)+~(C)*(~F*~E*D*B)*A+C*(~F*~E*D*B)*A)"),
    .INIT(64'hafafafafafaf27af))
    al_d848eac4 (
    .a(al_f5a4c6e6),
    .b(al_ee5ae3ff),
    .c(al_2802ceac),
    .d(al_a3de3eda[0]),
    .e(al_a3de3eda[2]),
    .f(al_a3de3eda[3]),
    .o(al_45c565e6));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(F)*~((~E*D*~C*~B))+~A*F*~((~E*D*~C*~B))+~(~A)*F*(~E*D*~C*~B)+~A*F*(~E*D*~C*~B))"),
    .INIT(64'h5555575555555455))
    al_ca59c0be (
    .a(al_45c565e6),
    .b(al_549b2fd9[0]),
    .c(al_549b2fd9[1]),
    .d(al_549b2fd9[2]),
    .e(al_549b2fd9[3]),
    .f(al_a6bbd516[0]),
    .o(al_fa675d9c));
  AL_DFF_X al_c00c07e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_fbb53e44),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a45b58d1));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(~C*B))"),
    .INIT(8'hae))
    al_b87f6b99 (
    .a(al_18c565c8),
    .b(al_a45b58d1),
    .c(al_e7b5abb5),
    .o(al_fbb53e44));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_96eb9d2c (
    .a(al_3d334d88),
    .b(al_36a894af[7]),
    .o(al_cac83419[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f1eee870 (
    .a(al_3d334d88),
    .b(al_36a894af[8]),
    .o(al_cac83419[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_24bc038c (
    .a(al_3d334d88),
    .b(al_36a894af[9]),
    .o(al_cac83419[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_9c2a79a7 (
    .a(al_3d334d88),
    .b(al_36a894af[10]),
    .o(al_cac83419[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_de92e263 (
    .a(al_3d334d88),
    .b(al_36a894af[11]),
    .o(al_cac83419[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_49124d1e (
    .a(al_6fd79ca[0]),
    .b(al_3d334d88),
    .o(al_63edc714[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_20a59860 (
    .a(al_6fd79ca[10]),
    .b(al_3d334d88),
    .o(al_63edc714[10]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_912710a1 (
    .a(al_6fd79ca[11]),
    .b(al_3d334d88),
    .o(al_63edc714[11]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_32337f5f (
    .a(al_6fd79ca[12]),
    .b(al_3d334d88),
    .o(al_63edc714[12]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_86fba2b6 (
    .a(al_6fd79ca[13]),
    .b(al_3d334d88),
    .o(al_63edc714[13]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_74796f33 (
    .a(al_6fd79ca[14]),
    .b(al_3d334d88),
    .o(al_63edc714[14]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_d30c5e1d (
    .a(al_6fd79ca[15]),
    .b(al_3d334d88),
    .o(al_63edc714[15]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_abca7107 (
    .a(al_6fd79ca[16]),
    .b(al_3d334d88),
    .o(al_63edc714[16]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_25fdc52e (
    .a(al_6fd79ca[17]),
    .b(al_3d334d88),
    .o(al_63edc714[17]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_af8c3f06 (
    .a(al_6fd79ca[18]),
    .b(al_3d334d88),
    .o(al_63edc714[18]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_a302126e (
    .a(al_6fd79ca[19]),
    .b(al_3d334d88),
    .o(al_63edc714[19]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_237fbc24 (
    .a(al_6fd79ca[1]),
    .b(al_3d334d88),
    .o(al_63edc714[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_7d6c5614 (
    .a(al_6fd79ca[20]),
    .b(al_3d334d88),
    .o(al_63edc714[20]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_c40d44e8 (
    .a(al_6fd79ca[21]),
    .b(al_3d334d88),
    .o(al_63edc714[21]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_7116b3d3 (
    .a(al_6fd79ca[22]),
    .b(al_3d334d88),
    .o(al_63edc714[22]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_1b6a2d1b (
    .a(al_6fd79ca[23]),
    .b(al_3d334d88),
    .o(al_63edc714[23]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_c7dc5297 (
    .a(al_6fd79ca[24]),
    .b(al_3d334d88),
    .o(al_63edc714[24]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_b3da0ad4 (
    .a(al_6fd79ca[25]),
    .b(al_3d334d88),
    .o(al_63edc714[25]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_88c3d2e5 (
    .a(al_6fd79ca[26]),
    .b(al_3d334d88),
    .o(al_63edc714[26]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_98ea21ea (
    .a(al_6fd79ca[27]),
    .b(al_3d334d88),
    .o(al_63edc714[27]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_aa4584b (
    .a(al_6fd79ca[28]),
    .b(al_3d334d88),
    .o(al_63edc714[28]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_be8647fa (
    .a(al_6fd79ca[29]),
    .b(al_3d334d88),
    .o(al_63edc714[29]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_a0e6539a (
    .a(al_6fd79ca[2]),
    .b(al_3d334d88),
    .o(al_63edc714[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_89372389 (
    .a(al_6fd79ca[30]),
    .b(al_3d334d88),
    .o(al_63edc714[30]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_c059744c (
    .a(al_6fd79ca[31]),
    .b(al_3d334d88),
    .o(al_63edc714[31]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_f3b8f310 (
    .a(al_6fd79ca[3]),
    .b(al_3d334d88),
    .o(al_63edc714[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_4d10718e (
    .a(al_6fd79ca[4]),
    .b(al_3d334d88),
    .o(al_63edc714[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_3fe5800d (
    .a(al_6fd79ca[5]),
    .b(al_3d334d88),
    .o(al_63edc714[5]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_cc1e2b0b (
    .a(al_6fd79ca[6]),
    .b(al_3d334d88),
    .o(al_63edc714[6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_73d516fb (
    .a(al_6fd79ca[7]),
    .b(al_3d334d88),
    .o(al_63edc714[7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_ed666f24 (
    .a(al_6fd79ca[8]),
    .b(al_3d334d88),
    .o(al_63edc714[8]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_724c1e45 (
    .a(al_6fd79ca[9]),
    .b(al_3d334d88),
    .o(al_63edc714[9]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_c954b48a (
    .a(al_5493f072),
    .b(al_3d334d88),
    .o(al_f36bf4fd));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*B*~(C)+A*B*~(C)+A*~(B)*C)"),
    .INIT(8'h2c))
    al_bf4bfaad (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_1d392f4f[0]),
    .o(al_2d4f70b0[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0afa3000))
    al_2b76ecc7 (
    .a(al_1d840c32),
    .b(al_cb40733a),
    .c(al_a430e4d2),
    .d(al_1d392f4f[0]),
    .e(al_1d392f4f[1]),
    .o(al_2d4f70b0[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h2ec0))
    al_e0697d50 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_92bdd050),
    .d(al_1d392f4f[2]),
    .o(al_2d4f70b0[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*(D*C)*~(E)+A*B*(D*C)*~(E)+A*~(B)*~((D*C))*E+~(A)*B*~((D*C))*E+A*B*~((D*C))*E+A*~(B)*(D*C)*E)"),
    .INIT(32'h2eeec000))
    al_653a9556 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_92bdd050),
    .d(al_1d392f4f[2]),
    .e(al_1d392f4f[3]),
    .o(al_2d4f70b0[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*(E*D*C)*~(F)+A*B*(E*D*C)*~(F)+A*~(B)*~((E*D*C))*F+~(A)*B*~((E*D*C))*F+A*B*~((E*D*C))*F+A*~(B)*(E*D*C)*F)"),
    .INIT(64'h2eeeeeeec0000000))
    al_720a3164 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_92bdd050),
    .d(al_1d392f4f[2]),
    .e(al_1d392f4f[3]),
    .f(al_1d392f4f[4]),
    .o(al_2d4f70b0[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_80537a55 (
    .a(al_1d392f4f[0]),
    .b(al_1d392f4f[1]),
    .o(al_92bdd050));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    al_f52321c4 (
    .a(al_1d392f4f[1]),
    .b(al_1d392f4f[2]),
    .c(al_1d392f4f[3]),
    .d(al_1d392f4f[4]),
    .e(al_1d392f4f[5]),
    .o(al_cb40733a));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_69c44458 (
    .a(al_a430e4d2),
    .b(al_92bdd050),
    .c(al_1d392f4f[2]),
    .d(al_1d392f4f[3]),
    .e(al_1d392f4f[4]),
    .o(al_4348da93));
  AL_MAP_LUT6 #(
    .EQN("(~(~B*~((E*C))*~(D)+~B*(E*C)*~(D)+~(~B)*(E*C)*D+~B*(E*C)*D)*(F@A))"),
    .INIT(64'h054455440a88aa88))
    al_1a7e2775 (
    .a(al_4348da93),
    .b(al_1d840c32),
    .c(al_cb40733a),
    .d(al_a430e4d2),
    .e(al_1d392f4f[0]),
    .f(al_1d392f4f[5]),
    .o(al_2d4f70b0[5]));
  AL_DFF_X al_8ddc2e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9cf531f8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9526c852));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    al_8b0214be (
    .a(al_bb0cd305),
    .b(al_6c5ae138),
    .c(al_9526c852),
    .o(al_9cf531f8));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_5c37af93 (
    .a(al_3e46fbe7),
    .b(al_60dd36d7),
    .o(al_ba08f61a));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_fd71327 (
    .a(al_3ebb68c3),
    .b(al_98804c07),
    .c(al_6d92b3c6),
    .d(al_bdb28b76),
    .e(al_73fb1ee5),
    .f(al_33a2911e),
    .o(al_eddc4d82));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_48f43cd9 (
    .a(al_d76255c5),
    .b(al_7d27d680),
    .c(al_f61ec828),
    .d(al_7e6320f4),
    .e(al_e6455839),
    .f(al_d00a6f56),
    .o(al_84c23d54));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_5a76fcb8 (
    .a(al_62da7380),
    .b(al_524d11ae),
    .c(al_eddc4d82),
    .d(al_84c23d54),
    .o(al_b968fef9));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B@(~D*C)))"),
    .INIT(16'h4414))
    al_5de192c9 (
    .a(al_b968fef9),
    .b(al_698ba8c2),
    .c(al_ba08f61a),
    .d(dBusAhb_HSIZE[1]),
    .o(al_86466d94));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_5ffc1a26 (
    .a(al_c5b8f9ea),
    .b(al_3e46fbe7),
    .c(al_14b732b9),
    .o(al_698ba8c2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_950ad2c (
    .a(al_1f5093b5),
    .b(al_ffc4fe26),
    .c(al_658bb789),
    .d(al_a831c176),
    .e(al_c7df4b4d),
    .f(al_3b0f4da7),
    .o(al_76ffd29c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_eb2c001e (
    .a(al_3626cb0),
    .b(al_3b8c31d7),
    .c(al_102b7ad2),
    .d(al_6ec45564),
    .e(al_e611ec68),
    .f(al_53b3dbc6),
    .o(al_def94157));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_6c271891 (
    .a(al_76ffd29c),
    .b(al_def94157),
    .c(dBusAhb_HSIZE[1]),
    .d(al_60dd36d7),
    .e(al_f1bb92e9),
    .o(al_62da7380));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_25cbef57 (
    .a(al_8a841cb4),
    .b(al_c861c8f0),
    .c(al_76a52f3d),
    .d(al_bf952132),
    .e(al_2370214),
    .f(al_f4b5275b),
    .o(al_524d11ae));
  AL_DFF_X al_8cb5138d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_86466d94),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a167c8cf));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_313264c2 (
    .a(al_b70cb9be[31]),
    .b(al_a5f7e6c[0]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b15a1641 (
    .a(al_7b59c46e[9]),
    .b(al_a5f7e6c[10]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8dfc7427 (
    .a(al_7b59c46e[10]),
    .b(al_a5f7e6c[11]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_91888681 (
    .a(al_7b59c46e[11]),
    .b(al_a5f7e6c[12]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4e2dcae3 (
    .a(al_7b59c46e[12]),
    .b(al_a5f7e6c[13]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d1dd8e2d (
    .a(al_7b59c46e[13]),
    .b(al_a5f7e6c[14]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_aa0b8e5d (
    .a(al_7b59c46e[14]),
    .b(al_a5f7e6c[15]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d34cb63 (
    .a(al_7b59c46e[15]),
    .b(al_a5f7e6c[16]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_53054297 (
    .a(al_7b59c46e[16]),
    .b(al_a5f7e6c[17]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_d2d40886 (
    .a(al_7b59c46e[17]),
    .b(al_a5f7e6c[18]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7621adaf (
    .a(al_7b59c46e[18]),
    .b(al_a5f7e6c[19]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e108040f (
    .a(al_7b59c46e[0]),
    .b(al_a5f7e6c[1]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a4a23576 (
    .a(al_7b59c46e[19]),
    .b(al_a5f7e6c[20]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5542d006 (
    .a(al_7b59c46e[20]),
    .b(al_a5f7e6c[21]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_2210c845 (
    .a(al_7b59c46e[21]),
    .b(al_a5f7e6c[22]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_6a005d44 (
    .a(al_7b59c46e[22]),
    .b(al_a5f7e6c[23]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5ee6f219 (
    .a(al_7b59c46e[23]),
    .b(al_a5f7e6c[24]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_91fe2d21 (
    .a(al_7b59c46e[24]),
    .b(al_a5f7e6c[25]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8d1b270a (
    .a(al_7b59c46e[25]),
    .b(al_a5f7e6c[26]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5fbd8b7b (
    .a(al_7b59c46e[26]),
    .b(al_a5f7e6c[27]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_c4b1eb92 (
    .a(al_7b59c46e[27]),
    .b(al_a5f7e6c[28]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_6168e814 (
    .a(al_7b59c46e[28]),
    .b(al_a5f7e6c[29]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_753dc118 (
    .a(al_7b59c46e[1]),
    .b(al_a5f7e6c[2]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_188fdbb5 (
    .a(al_7b59c46e[29]),
    .b(al_a5f7e6c[30]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_8911aab4 (
    .a(al_7b59c46e[30]),
    .b(al_a5f7e6c[31]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a599bf39 (
    .a(al_7b59c46e[2]),
    .b(al_a5f7e6c[3]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b0cf0be (
    .a(al_7b59c46e[3]),
    .b(al_a5f7e6c[4]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5e71bdfa (
    .a(al_7b59c46e[4]),
    .b(al_a5f7e6c[5]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_557507b9 (
    .a(al_7b59c46e[5]),
    .b(al_a5f7e6c[6]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_42b022d8 (
    .a(al_7b59c46e[6]),
    .b(al_a5f7e6c[7]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_cc0a43e4 (
    .a(al_7b59c46e[7]),
    .b(al_a5f7e6c[8]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_284a4531 (
    .a(al_7b59c46e[8]),
    .b(al_a5f7e6c[9]),
    .c(al_a5f7e6c[32]),
    .o(al_830b3656[9]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_6a0540d4 (
    .a(al_698ba8c2),
    .b(al_1891b3c7),
    .o(al_439698e9[0]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_6245ec1b (
    .a(al_698ba8c2),
    .b(al_407c8ac1),
    .o(al_439698e9[10]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_7a6f64cf (
    .a(al_698ba8c2),
    .b(al_fdf9f0dc),
    .o(al_439698e9[11]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_879999ff (
    .a(al_698ba8c2),
    .b(al_b5bf2603),
    .o(al_439698e9[12]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_d5b342c1 (
    .a(al_698ba8c2),
    .b(al_c8ba6c61),
    .o(al_439698e9[13]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_4a394eee (
    .a(al_698ba8c2),
    .b(al_59be2ab1),
    .o(al_439698e9[14]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_2ac75922 (
    .a(al_698ba8c2),
    .b(al_8488923),
    .o(al_439698e9[15]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_bbf19c78 (
    .a(al_698ba8c2),
    .b(al_5727b773),
    .o(al_439698e9[16]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_4d0644a2 (
    .a(al_698ba8c2),
    .b(al_eead7739),
    .o(al_439698e9[17]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_c1ec2522 (
    .a(al_698ba8c2),
    .b(al_f430a5aa),
    .o(al_439698e9[18]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_1ed460b6 (
    .a(al_698ba8c2),
    .b(al_cd498e9f),
    .o(al_439698e9[19]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_60cf99be (
    .a(al_698ba8c2),
    .b(al_512b1421),
    .o(al_439698e9[1]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e89f90aa (
    .a(al_698ba8c2),
    .b(al_3656d228),
    .o(al_439698e9[20]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_96a15db7 (
    .a(al_698ba8c2),
    .b(al_30f08f9c),
    .o(al_439698e9[21]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_1728eac (
    .a(al_698ba8c2),
    .b(al_bf6a3977),
    .o(al_439698e9[22]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_5e870b02 (
    .a(al_698ba8c2),
    .b(al_2ede456b),
    .o(al_439698e9[23]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_99addeda (
    .a(al_698ba8c2),
    .b(al_3a7c5a5),
    .o(al_439698e9[24]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_ac0cd29d (
    .a(al_698ba8c2),
    .b(al_9b707062),
    .o(al_439698e9[25]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_7d750fec (
    .a(al_698ba8c2),
    .b(al_a69cec28),
    .o(al_439698e9[26]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_863bd294 (
    .a(al_698ba8c2),
    .b(al_d78f6bd4),
    .o(al_439698e9[27]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_3caa0801 (
    .a(al_698ba8c2),
    .b(al_cae21d2e),
    .o(al_439698e9[28]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_ec7fa1d5 (
    .a(al_698ba8c2),
    .b(al_19c0990d),
    .o(al_439698e9[29]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_1e1650f (
    .a(al_698ba8c2),
    .b(al_80e2c141),
    .o(al_439698e9[2]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e9f35bf2 (
    .a(al_698ba8c2),
    .b(al_cacb44c4),
    .o(al_439698e9[30]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_7c4e046b (
    .a(al_698ba8c2),
    .b(al_14b732b9),
    .o(al_439698e9[31]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_fff9b3dc (
    .a(al_698ba8c2),
    .b(al_1e979a01),
    .o(al_439698e9[3]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_17ae26dc (
    .a(al_698ba8c2),
    .b(al_5df930ee),
    .o(al_439698e9[4]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_ef770a75 (
    .a(al_698ba8c2),
    .b(al_8e267e24),
    .o(al_439698e9[5]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_25c44dd1 (
    .a(al_698ba8c2),
    .b(al_e163f204),
    .o(al_439698e9[6]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_d295fb9 (
    .a(al_698ba8c2),
    .b(al_a6e0ed04),
    .o(al_439698e9[7]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_d8e6d3dc (
    .a(al_698ba8c2),
    .b(al_a35cf148),
    .o(al_439698e9[8]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_230296b0 (
    .a(al_698ba8c2),
    .b(al_728c73ac),
    .o(al_439698e9[9]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(C)*~(A)+E*C*~(A)+~(E)*C*A+E*C*A)*~(D)*~(B)+~(E*~(C)*~(A)+E*C*~(A)+~(E)*C*A+E*C*A)*D*~(B)+~(~(E*~(C)*~(A)+E*C*~(A)+~(E)*C*A+E*C*A))*D*B+~(E*~(C)*~(A)+E*C*~(A)+~(E)*C*A+E*C*A)*D*B)"),
    .INIT(32'h31fd20ec))
    al_675f4059 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_b70cb9be[0]),
    .d(al_a5f7e6c[32]),
    .e(al_1891b3c7),
    .o(al_d0c02c51[0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_26ca761e (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[10]),
    .d(al_b70cb9be[9]),
    .e(al_b70cb9be[10]),
    .o(al_d0c02c51[10]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_4ba9c671 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[11]),
    .d(al_b70cb9be[10]),
    .e(al_b70cb9be[11]),
    .o(al_d0c02c51[11]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_c13a0934 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[12]),
    .d(al_b70cb9be[11]),
    .e(al_b70cb9be[12]),
    .o(al_d0c02c51[12]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_e93cfc02 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[13]),
    .d(al_b70cb9be[12]),
    .e(al_b70cb9be[13]),
    .o(al_d0c02c51[13]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_b41e171e (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[14]),
    .d(al_b70cb9be[13]),
    .e(al_b70cb9be[14]),
    .o(al_d0c02c51[14]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_724bfc94 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[15]),
    .d(al_b70cb9be[14]),
    .e(al_b70cb9be[15]),
    .o(al_d0c02c51[15]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_11d3a0eb (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[16]),
    .d(al_b70cb9be[15]),
    .e(al_b70cb9be[16]),
    .o(al_d0c02c51[16]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_2683c6b9 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[17]),
    .d(al_b70cb9be[16]),
    .e(al_b70cb9be[17]),
    .o(al_d0c02c51[17]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_e557a608 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[18]),
    .d(al_b70cb9be[17]),
    .e(al_b70cb9be[18]),
    .o(al_d0c02c51[18]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_a3c2e5b8 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[19]),
    .d(al_b70cb9be[18]),
    .e(al_b70cb9be[19]),
    .o(al_d0c02c51[19]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_8d42411a (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[1]),
    .d(al_b70cb9be[0]),
    .e(al_b70cb9be[1]),
    .o(al_d0c02c51[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_b5a2ecf2 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[20]),
    .d(al_b70cb9be[19]),
    .e(al_b70cb9be[20]),
    .o(al_d0c02c51[20]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_7e739d4d (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[21]),
    .d(al_b70cb9be[20]),
    .e(al_b70cb9be[21]),
    .o(al_d0c02c51[21]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_eb9a8768 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[22]),
    .d(al_b70cb9be[21]),
    .e(al_b70cb9be[22]),
    .o(al_d0c02c51[22]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_eb2d7da3 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[23]),
    .d(al_b70cb9be[22]),
    .e(al_b70cb9be[23]),
    .o(al_d0c02c51[23]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_10960b6f (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[24]),
    .d(al_b70cb9be[23]),
    .e(al_b70cb9be[24]),
    .o(al_d0c02c51[24]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_930f88c0 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[25]),
    .d(al_b70cb9be[24]),
    .e(al_b70cb9be[25]),
    .o(al_d0c02c51[25]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_b2261a4e (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[26]),
    .d(al_b70cb9be[25]),
    .e(al_b70cb9be[26]),
    .o(al_d0c02c51[26]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_958dd28d (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[27]),
    .d(al_b70cb9be[26]),
    .e(al_b70cb9be[27]),
    .o(al_d0c02c51[27]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_ceccb84f (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[28]),
    .d(al_b70cb9be[27]),
    .e(al_b70cb9be[28]),
    .o(al_d0c02c51[28]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_e20f7942 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[29]),
    .d(al_b70cb9be[28]),
    .e(al_b70cb9be[29]),
    .o(al_d0c02c51[29]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_77176486 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[2]),
    .d(al_b70cb9be[1]),
    .e(al_b70cb9be[2]),
    .o(al_d0c02c51[2]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_2be1b21e (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[30]),
    .d(al_b70cb9be[29]),
    .e(al_b70cb9be[30]),
    .o(al_d0c02c51[30]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_82919e50 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[31]),
    .d(al_b70cb9be[30]),
    .e(al_b70cb9be[31]),
    .o(al_d0c02c51[31]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_5d5a9cff (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[3]),
    .d(al_b70cb9be[2]),
    .e(al_b70cb9be[3]),
    .o(al_d0c02c51[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_a552db15 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[4]),
    .d(al_b70cb9be[3]),
    .e(al_b70cb9be[4]),
    .o(al_d0c02c51[4]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_260a1ff4 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[5]),
    .d(al_b70cb9be[4]),
    .e(al_b70cb9be[5]),
    .o(al_d0c02c51[5]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_da2bb8bf (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[6]),
    .d(al_b70cb9be[5]),
    .e(al_b70cb9be[6]),
    .o(al_d0c02c51[6]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_11679f4 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[7]),
    .d(al_b70cb9be[6]),
    .e(al_b70cb9be[7]),
    .o(al_d0c02c51[7]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_61a0a172 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[8]),
    .d(al_b70cb9be[7]),
    .e(al_b70cb9be[8]),
    .o(al_d0c02c51[8]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(D)*~(B)+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*~(B)+~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*D*B+(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*D*B)"),
    .INIT(32'hfe32dc10))
    al_56da65a4 (
    .a(al_1d840c32),
    .b(al_a430e4d2),
    .c(al_afda7fe3[9]),
    .d(al_b70cb9be[8]),
    .e(al_b70cb9be[9]),
    .o(al_d0c02c51[9]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_4e6e1793 (
    .a(al_ba08f61a),
    .b(al_f4b5275b),
    .o(al_4e7a070d[0]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_56416670 (
    .a(al_ba08f61a),
    .b(al_98804c07),
    .o(al_4e7a070d[10]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_d96a064f (
    .a(al_ba08f61a),
    .b(al_3ebb68c3),
    .o(al_4e7a070d[11]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_1da07387 (
    .a(al_ba08f61a),
    .b(al_d00a6f56),
    .o(al_4e7a070d[12]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_c718e7aa (
    .a(al_ba08f61a),
    .b(al_e6455839),
    .o(al_4e7a070d[13]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_230e8e37 (
    .a(al_ba08f61a),
    .b(al_7e6320f4),
    .o(al_4e7a070d[14]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e2841ae4 (
    .a(al_ba08f61a),
    .b(al_f61ec828),
    .o(al_4e7a070d[15]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_674967df (
    .a(al_ba08f61a),
    .b(al_7d27d680),
    .o(al_4e7a070d[16]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_258290ec (
    .a(al_ba08f61a),
    .b(al_d76255c5),
    .o(al_4e7a070d[17]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_68707dd4 (
    .a(al_ba08f61a),
    .b(al_3b0f4da7),
    .o(al_4e7a070d[18]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_5cb31166 (
    .a(al_ba08f61a),
    .b(al_c7df4b4d),
    .o(al_4e7a070d[19]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_5f3632c1 (
    .a(al_ba08f61a),
    .b(al_2370214),
    .o(al_4e7a070d[1]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_c555e9d3 (
    .a(al_ba08f61a),
    .b(al_a831c176),
    .o(al_4e7a070d[20]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_380117e1 (
    .a(al_ba08f61a),
    .b(al_658bb789),
    .o(al_4e7a070d[21]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_2e8c4a9d (
    .a(al_ba08f61a),
    .b(al_ffc4fe26),
    .o(al_4e7a070d[22]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_a36922b6 (
    .a(al_ba08f61a),
    .b(al_1f5093b5),
    .o(al_4e7a070d[23]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_acc7f5ea (
    .a(al_ba08f61a),
    .b(al_53b3dbc6),
    .o(al_4e7a070d[24]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_2e1ce069 (
    .a(al_ba08f61a),
    .b(al_e611ec68),
    .o(al_4e7a070d[25]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_bf7bc2bb (
    .a(al_ba08f61a),
    .b(al_6ec45564),
    .o(al_4e7a070d[26]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_7742a418 (
    .a(al_ba08f61a),
    .b(al_102b7ad2),
    .o(al_4e7a070d[27]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_763b0177 (
    .a(al_ba08f61a),
    .b(al_3b8c31d7),
    .o(al_4e7a070d[28]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_66a404d2 (
    .a(al_ba08f61a),
    .b(al_3626cb0),
    .o(al_4e7a070d[29]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_2301f7d0 (
    .a(al_ba08f61a),
    .b(al_bf952132),
    .o(al_4e7a070d[2]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_32b65261 (
    .a(al_ba08f61a),
    .b(al_f1bb92e9),
    .o(al_4e7a070d[30]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e868150f (
    .a(al_3e46fbe7),
    .b(al_60dd36d7),
    .o(al_4e7a070d[31]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_ff972a8 (
    .a(al_ba08f61a),
    .b(al_76a52f3d),
    .o(al_4e7a070d[3]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_94b89bf9 (
    .a(al_ba08f61a),
    .b(al_c861c8f0),
    .o(al_4e7a070d[4]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_d8278efd (
    .a(al_ba08f61a),
    .b(al_8a841cb4),
    .o(al_4e7a070d[5]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_65a30f8e (
    .a(al_ba08f61a),
    .b(al_33a2911e),
    .o(al_4e7a070d[6]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_7e593d96 (
    .a(al_ba08f61a),
    .b(al_73fb1ee5),
    .o(al_4e7a070d[7]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_a2630eb2 (
    .a(al_ba08f61a),
    .b(al_bdb28b76),
    .o(al_4e7a070d[8]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_bf3a386a (
    .a(al_ba08f61a),
    .b(al_6d92b3c6),
    .o(al_4e7a070d[9]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_95eb934a (
    .a(al_bb0cd305),
    .o(al_98842338));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*C*B)*~(~D*A))"),
    .INIT(32'hc0ea00aa))
    al_9ee79242 (
    .a(al_1a1af7e4),
    .b(al_592c9a6),
    .c(al_5a744f0f),
    .d(al_bb0cd305),
    .e(al_523cde28),
    .o(al_82faef35));
  AL_DFF_X al_9dc100f3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_82faef35),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_501dbbdf));
  AL_DFF_X al_1618478b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e3290619),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41e75372));
  AL_DFF_X al_96366f5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e3edcf1a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2af4b91));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_8de01616 (
    .a(1'b0),
    .o({al_428c2665,open_n47}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7b9ad123 (
    .a(al_1d8f7667[0]),
    .b(al_71c7f8f0[32]),
    .c(al_428c2665),
    .o({al_77af043a,al_d7ecfd18[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8d97dc59 (
    .a(al_1d8f7667[1]),
    .b(al_71c7f8f0[33]),
    .c(al_77af043a),
    .o({al_c99791ac,al_d7ecfd18[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_62530da0 (
    .a(al_1d8f7667[2]),
    .b(al_71c7f8f0[34]),
    .c(al_c99791ac),
    .o({al_18a866ae,al_d7ecfd18[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_82283be1 (
    .a(al_1d8f7667[3]),
    .b(al_71c7f8f0[35]),
    .c(al_18a866ae),
    .o({al_9cb94e30,al_d7ecfd18[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_666d0567 (
    .a(al_1d8f7667[4]),
    .b(al_71c7f8f0[36]),
    .c(al_9cb94e30),
    .o({al_1e7370cf,al_d7ecfd18[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4ca40e36 (
    .a(al_1d8f7667[5]),
    .b(al_71c7f8f0[37]),
    .c(al_1e7370cf),
    .o({al_1712bb7c,al_d7ecfd18[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_30aa2e88 (
    .a(al_1d8f7667[6]),
    .b(al_71c7f8f0[38]),
    .c(al_1712bb7c),
    .o({al_3043d922,al_d7ecfd18[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c2e81cdc (
    .a(al_1d8f7667[7]),
    .b(al_71c7f8f0[39]),
    .c(al_3043d922),
    .o({al_69790d6e,al_d7ecfd18[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fd4e6cb0 (
    .a(al_1d8f7667[8]),
    .b(al_71c7f8f0[40]),
    .c(al_69790d6e),
    .o({al_b1c0d1f7,al_d7ecfd18[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4b929999 (
    .a(al_1d8f7667[9]),
    .b(al_71c7f8f0[41]),
    .c(al_b1c0d1f7),
    .o({al_58533fed,al_d7ecfd18[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_91a7faa2 (
    .a(al_1d8f7667[10]),
    .b(al_71c7f8f0[42]),
    .c(al_58533fed),
    .o({al_fa53107d,al_d7ecfd18[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e7581646 (
    .a(al_1d8f7667[11]),
    .b(al_71c7f8f0[43]),
    .c(al_fa53107d),
    .o({al_7a87cf81,al_d7ecfd18[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bb0de5c2 (
    .a(al_1d8f7667[12]),
    .b(al_71c7f8f0[44]),
    .c(al_7a87cf81),
    .o({al_3ca77acd,al_d7ecfd18[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_589babdd (
    .a(al_1d8f7667[13]),
    .b(al_71c7f8f0[45]),
    .c(al_3ca77acd),
    .o({al_19663434,al_d7ecfd18[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e6430f30 (
    .a(al_1d8f7667[14]),
    .b(al_71c7f8f0[46]),
    .c(al_19663434),
    .o({al_8e3e7ef7,al_d7ecfd18[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6a92233b (
    .a(al_1d8f7667[15]),
    .b(al_71c7f8f0[47]),
    .c(al_8e3e7ef7),
    .o({al_1df72327,al_d7ecfd18[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_538f8ff6 (
    .a(al_1d8f7667[16]),
    .b(al_71c7f8f0[48]),
    .c(al_1df72327),
    .o({al_f07170fc,al_d7ecfd18[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bfd2edc0 (
    .a(al_1d8f7667[17]),
    .b(al_71c7f8f0[49]),
    .c(al_f07170fc),
    .o({al_5632987e,al_d7ecfd18[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_937e6e92 (
    .a(al_1d8f7667[18]),
    .b(al_71c7f8f0[50]),
    .c(al_5632987e),
    .o({al_c5c038e7,al_d7ecfd18[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1af27a78 (
    .a(al_1d8f7667[19]),
    .b(al_71c7f8f0[51]),
    .c(al_c5c038e7),
    .o({al_e56ae954,al_d7ecfd18[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b2c4716e (
    .a(al_1d8f7667[20]),
    .b(al_71c7f8f0[51]),
    .c(al_e56ae954),
    .o({al_83a5fe89,al_d7ecfd18[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_59390ce (
    .a(al_1d8f7667[21]),
    .b(al_71c7f8f0[51]),
    .c(al_83a5fe89),
    .o({al_ad72d731,al_d7ecfd18[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3cd9ce70 (
    .a(al_1d8f7667[22]),
    .b(al_71c7f8f0[51]),
    .c(al_ad72d731),
    .o({al_e6ba0c27,al_d7ecfd18[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_88e686cb (
    .a(al_1d8f7667[23]),
    .b(al_71c7f8f0[51]),
    .c(al_e6ba0c27),
    .o({al_41cca93a,al_d7ecfd18[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_729b5703 (
    .a(al_1d8f7667[24]),
    .b(al_71c7f8f0[51]),
    .c(al_41cca93a),
    .o({al_19790099,al_d7ecfd18[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3ae513d6 (
    .a(al_1d8f7667[25]),
    .b(al_71c7f8f0[51]),
    .c(al_19790099),
    .o({al_ab63694b,al_d7ecfd18[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f42a56d6 (
    .a(al_1d8f7667[26]),
    .b(al_71c7f8f0[51]),
    .c(al_ab63694b),
    .o({al_35ca4317,al_d7ecfd18[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_75aa4a6e (
    .a(al_1d8f7667[27]),
    .b(al_71c7f8f0[51]),
    .c(al_35ca4317),
    .o({al_32a84555,al_d7ecfd18[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_226e4319 (
    .a(al_1d8f7667[28]),
    .b(al_71c7f8f0[51]),
    .c(al_32a84555),
    .o({al_9b78efe2,al_d7ecfd18[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ce0c3191 (
    .a(al_1d8f7667[29]),
    .b(al_71c7f8f0[51]),
    .c(al_9b78efe2),
    .o({al_4507eb5c,al_d7ecfd18[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7e81eadf (
    .a(al_1d8f7667[30]),
    .b(al_71c7f8f0[51]),
    .c(al_4507eb5c),
    .o({al_627e0d7d,al_d7ecfd18[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_86d674f8 (
    .a(al_1d8f7667[31]),
    .b(al_71c7f8f0[51]),
    .c(al_627e0d7d),
    .o({open_n48,al_d7ecfd18[31]}));
  AL_DFF_X al_807b8831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_24641d37),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca0e00e));
  PH1_PHY_DSPREG #(
    .CEMUX("INV"),
    .CLKMUX("SIG"),
    .RSTMODE("ASYNC"),
    .RSTMUX("0"),
    .WIDTH(45))
    al_d6352cbf (
    .ce(al_98842338),
    .clk(SYS_CLK),
    .d(al_de2ed994),
    .rst(1'bx),
    .q(al_9aa9386d));
  PH1_PHY_DSPREG #(
    .CEMUX("1"),
    .CLKMUX("SIG"),
    .RSTMODE("ASYNC"),
    .RSTMUX("0"),
    .WIDTH(54))
    al_27fd71f0 (
    .ce(1'bx),
    .clk(SYS_CLK),
    .d(al_25ac6d54),
    .rst(1'bx),
    .q({al_193295bb[53:32],al_1d8f7667[31:0]}));
  PH1_PHY_DSPMULT
    al_351527f9 (
    .opctrl(2'b11),
    .x({al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_14b732b9,al_cacb44c4,al_19c0990d,al_cae21d2e,al_d78f6bd4,al_a69cec28,al_9b707062,al_3a7c5a5,al_2ede456b,al_bf6a3977,al_30f08f9c,al_3656d228,al_cd498e9f,al_f430a5aa,al_eead7739,al_5727b773}),
    .y({al_65e3dd93[16],al_65e3dd93[16],al_60dd36d7,al_f1bb92e9,al_3626cb0,al_3b8c31d7,al_102b7ad2,al_6ec45564,al_e611ec68,al_53b3dbc6,al_1f5093b5,al_ffc4fe26,al_658bb789,al_a831c176,al_c7df4b4d,al_3b0f4da7,al_d76255c5,al_7d27d680}),
    .p(al_de2ed994));
  PH1_PHY_DSPTADD #(
    .CI_INVERT("NO"),
    .INV_OPCTRL(4'b0000),
    .RND_CONST(54'b0),
    .USE_OVERFLOW("S53"),
    .X1_EXTEND("YES"),
    .Y1_ROUND("NO"),
    .Z1_SHIFT("NO"))
    al_b64c0b48 (
    .ci(1'b0),
    .ci_special(1'b0),
    .opctrl(9'b000100000),
    .x1_special({al_9aa9386d[44],al_9aa9386d[44],al_9aa9386d[44],al_9aa9386d[44],al_9aa9386d[44],al_9aa9386d[44],al_9aa9386d[44],al_9aa9386d[44],al_9aa9386d[44],al_9aa9386d}),
    .y0(54'b000000000000000000000000000000000000000000000000000000),
    .y1_special(54'b000000000000000000000000000000000000000000000000000000),
    .z0(54'b000000000000000000000000000000000000000000000000000000),
    .z1_special(54'b000000000000000000000000000000000000000000000000000000),
    .sum(al_25ac6d54));
  PH1_PHY_DSPREG #(
    .CEMUX("INV"),
    .CLKMUX("SIG"),
    .RSTMODE("ASYNC"),
    .RSTMUX("0"),
    .WIDTH(45))
    al_32773bd8 (
    .ce(al_98842338),
    .clk(SYS_CLK),
    .d(al_1ee074c7),
    .rst(1'bx),
    .q({al_63395efb[44:34],al_3d2fbc2e}));
  PH1_PHY_DSPMULT
    al_ef007631 (
    .opctrl(2'b11),
    .x({al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_da34572b[16],al_14b732b9,al_cacb44c4,al_19c0990d,al_cae21d2e,al_d78f6bd4,al_a69cec28,al_9b707062,al_3a7c5a5,al_2ede456b,al_bf6a3977,al_30f08f9c,al_3656d228,al_cd498e9f,al_f430a5aa,al_eead7739,al_5727b773}),
    .y({2'b00,al_f61ec828,al_7e6320f4,al_e6455839,al_d00a6f56,al_3ebb68c3,al_98804c07,al_6d92b3c6,al_bdb28b76,al_73fb1ee5,al_33a2911e,al_8a841cb4,al_c861c8f0,al_76a52f3d,al_bf952132,al_2370214,al_f4b5275b}),
    .p(al_1ee074c7));
  PH1_PHY_DSPREG #(
    .CEMUX("INV"),
    .CLKMUX("SIG"),
    .RSTMODE("ASYNC"),
    .RSTMUX("0"),
    .WIDTH(45))
    al_e40ca92a (
    .ce(al_98842338),
    .clk(SYS_CLK),
    .d(al_8ffa2af5),
    .rst(1'bx),
    .q({al_186e4c3b[44:34],al_9edb1d1e}));
  PH1_PHY_DSPMULT
    al_2e57b26 (
    .opctrl(2'b11),
    .x({11'b00000000000,al_8488923,al_59be2ab1,al_c8ba6c61,al_b5bf2603,al_fdf9f0dc,al_407c8ac1,al_728c73ac,al_a35cf148,al_a6e0ed04,al_e163f204,al_8e267e24,al_5df930ee,al_1e979a01,al_80e2c141,al_512b1421,al_1891b3c7}),
    .y({al_65e3dd93[16],al_65e3dd93[16],al_60dd36d7,al_f1bb92e9,al_3626cb0,al_3b8c31d7,al_102b7ad2,al_6ec45564,al_e611ec68,al_53b3dbc6,al_1f5093b5,al_ffc4fe26,al_658bb789,al_a831c176,al_c7df4b4d,al_3b0f4da7,al_d76255c5,al_7d27d680}),
    .p(al_8ffa2af5));
  PH1_PHY_DSPREG #(
    .CEMUX("INV"),
    .CLKMUX("SIG"),
    .RSTMODE("ASYNC"),
    .RSTMUX("0"),
    .WIDTH(45))
    al_cc5cb0ca (
    .ce(al_98842338),
    .clk(SYS_CLK),
    .d(al_3d954d6),
    .rst(1'bx),
    .q({al_4dc1fe7[44:32],al_ccb50b3a}));
  PH1_PHY_DSPMULT
    al_6a0906c8 (
    .opctrl(2'b11),
    .x({11'b00000000000,al_8488923,al_59be2ab1,al_c8ba6c61,al_b5bf2603,al_fdf9f0dc,al_407c8ac1,al_728c73ac,al_a35cf148,al_a6e0ed04,al_e163f204,al_8e267e24,al_5df930ee,al_1e979a01,al_80e2c141,al_512b1421,al_1891b3c7}),
    .y({2'b00,al_f61ec828,al_7e6320f4,al_e6455839,al_d00a6f56,al_3ebb68c3,al_98804c07,al_6d92b3c6,al_bdb28b76,al_73fb1ee5,al_33a2911e,al_8a841cb4,al_c861c8f0,al_76a52f3d,al_bf952132,al_2370214,al_f4b5275b}),
    .p(al_3d954d6));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_a749b0f8 (
    .a(al_9176d089),
    .b(al_d19b9f6b),
    .o(al_22883704));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_f82c2651 (
    .a(al_cb40733a),
    .b(al_1d392f4f[0]),
    .o(al_6c5ae138));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_c2373940 (
    .a(al_6c5ae138),
    .b(al_a430e4d2),
    .o(al_3f04848f));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(32),
    .DATA_WIDTH_W(32),
    .FILL_ALL("NONE"),
    .INIT_FILE("init_str:00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000"),
    .READREG("DISABLE"))
    al_3cb2d510 (
    .di(al_63edc714),
    .raddr(al_704d20e3[19:15]),
    .waddr(al_cac83419),
    .wclk(SYS_CLK),
    .we(al_f36bf4fd),
    .rdo(al_8c7f68e2));
  PH1_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(32),
    .DATA_WIDTH_W(32),
    .FILL_ALL("NONE"),
    .INIT_FILE("init_str:00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000 00000000000000000000000000000000"),
    .READREG("DISABLE"))
    al_d03d7d95 (
    .di(al_63edc714),
    .raddr(al_704d20e3[24:20]),
    .waddr(al_cac83419),
    .wclk(SYS_CLK),
    .we(al_f36bf4fd),
    .rdo(al_8492e16));
  AL_DFF_X al_cde7e75c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[8]));
  AL_DFF_X al_bcb8a13b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[9]));
  AL_DFF_X al_cf25ccc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[10]));
  AL_DFF_X al_3133f55f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[11]));
  AL_DFF_X al_6f36e1dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[12]));
  AL_DFF_X al_822a9ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[13]));
  AL_DFF_X al_b319db91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[14]));
  AL_DFF_X al_8ea71f14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[15]));
  AL_DFF_X al_5d315a33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[16]));
  AL_DFF_X al_38bf5476 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[17]));
  AL_DFF_X al_661193ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[0]));
  AL_DFF_X al_9437c821 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[18]));
  AL_DFF_X al_3194242c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[19]));
  AL_DFF_X al_d9587b8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[20]));
  AL_DFF_X al_8e638631 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[21]));
  AL_DFF_X al_9f8e7c72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[22]));
  AL_DFF_X al_cdd75e09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[23]));
  AL_DFF_X al_a1706ebe (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[24]));
  AL_DFF_X al_e0148ebe (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[25]));
  AL_DFF_X al_e0e496c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[26]));
  AL_DFF_X al_c2c5ad4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[27]));
  AL_DFF_X al_980c5972 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[1]));
  AL_DFF_X al_b8e0cf5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[28]));
  AL_DFF_X al_3ce6a918 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[29]));
  AL_DFF_X al_8a66cc42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[30]));
  AL_DFF_X al_e2c4f0cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[31]));
  AL_DFF_X al_a2a4fbfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[2]));
  AL_DFF_X al_859cf13a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[3]));
  AL_DFF_X al_686167be (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[4]));
  AL_DFF_X al_a1b48049 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[5]));
  AL_DFF_X al_9571a46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[6]));
  AL_DFF_X al_5b79bc56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3dcca8e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45e5d9f7[7]));
  AL_DFF_X al_ff304992 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[10]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[8]));
  AL_DFF_X al_1442714e (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[11]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[9]));
  AL_DFF_X al_e8034dc3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[12]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[10]));
  AL_DFF_X al_c7c31713 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[13]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[11]));
  AL_DFF_X al_3900d313 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[14]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[12]));
  AL_DFF_X al_908af27 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[15]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[13]));
  AL_DFF_X al_5246ea17 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[16]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[14]));
  AL_DFF_X al_d0114b25 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[17]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[15]));
  AL_DFF_X al_8b8c9274 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[18]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[16]));
  AL_DFF_X al_d56618c3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[19]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[17]));
  AL_DFF_X al_9dc3a88f (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[2]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[0]));
  AL_DFF_X al_cb6a5fc9 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[20]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[18]));
  AL_DFF_X al_d935accb (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[21]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[19]));
  AL_DFF_X al_5c85c5e6 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[22]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[20]));
  AL_DFF_X al_d569b387 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[23]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[21]));
  AL_DFF_X al_5a79cf86 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[24]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[22]));
  AL_DFF_X al_44b1cafd (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[25]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[23]));
  AL_DFF_X al_66fac08b (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[26]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[24]));
  AL_DFF_X al_1c328e59 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[27]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[25]));
  AL_DFF_X al_3ec74209 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[28]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[26]));
  AL_DFF_X al_a7f32229 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[29]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[27]));
  AL_DFF_X al_ad3c4ca8 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[3]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[1]));
  AL_DFF_X al_48f447ff (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[30]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[28]));
  AL_DFF_X al_2f82ce3e (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[31]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[29]));
  AL_DFF_X al_5cf2645f (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[4]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[2]));
  AL_DFF_X al_1d95c0a9 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[5]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[3]));
  AL_DFF_X al_3f4582a1 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[6]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[4]));
  AL_DFF_X al_f3cdbe6a (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[7]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[5]));
  AL_DFF_X al_49d30bfd (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[8]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[6]));
  AL_DFF_X al_b2fb79d6 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[9]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35d85285[7]));
  AL_DFF_X al_71dd1073 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[0]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41e76523[0]));
  AL_DFF_X al_a2f45ffa (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3bdbe1c8[1]),
    .en(al_22883704),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_41e76523[1]));
  AL_DFF_X al_93244f28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[8]));
  AL_DFF_X al_49918a9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[9]));
  AL_DFF_X al_d4adb855 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[10]));
  AL_DFF_X al_47d17b9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[11]));
  AL_DFF_X al_bd810d41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[12]));
  AL_DFF_X al_73759cf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[13]));
  AL_DFF_X al_e10d88a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[14]));
  AL_DFF_X al_501b9cc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[15]));
  AL_DFF_X al_17627450 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[16]));
  AL_DFF_X al_9193e662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[17]));
  AL_DFF_X al_9762ad7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[0]));
  AL_DFF_X al_1fa1d326 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[18]));
  AL_DFF_X al_4eb33c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[19]));
  AL_DFF_X al_92e22a21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[20]));
  AL_DFF_X al_ba24a737 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[21]));
  AL_DFF_X al_d0e611c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[22]));
  AL_DFF_X al_7b9f2b5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[23]));
  AL_DFF_X al_e817aaa8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[24]));
  AL_DFF_X al_46876c18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[25]));
  AL_DFF_X al_f289725d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[26]));
  AL_DFF_X al_7372d562 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[27]));
  AL_DFF_X al_b49534ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[1]));
  AL_DFF_X al_6661da7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[28]));
  AL_DFF_X al_661991aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[29]));
  AL_DFF_X al_3148a9eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[30]));
  AL_DFF_X al_a9071091 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[31]));
  AL_DFF_X al_f72b3b98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[2]));
  AL_DFF_X al_ad30cb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[3]));
  AL_DFF_X al_964d5e45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[4]));
  AL_DFF_X al_b9119904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[5]));
  AL_DFF_X al_6d941b44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[6]));
  AL_DFF_X al_164d0f2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d610ac57[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43722bf9[7]));
  AL_DFF_X al_2ffe404d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_36a894af[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a6a2b33[0]));
  AL_DFF_X al_fb048123 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_36a894af[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a6a2b33[1]));
  AL_DFF_X al_d48576a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_36a894af[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a6a2b33[2]));
  AL_DFF_X al_e1954430 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_36a894af[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a6a2b33[3]));
  AL_DFF_X al_d5b136f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_36a894af[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a6a2b33[4]));
  AL_DFF_X al_f99831ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[8]));
  AL_DFF_X al_35e6bab3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[9]));
  AL_DFF_X al_319233f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[10]));
  AL_DFF_X al_cb8264a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[11]));
  AL_DFF_X al_55db45b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[12]));
  AL_DFF_X al_42a068c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[13]));
  AL_DFF_X al_ce680d74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[14]));
  AL_DFF_X al_5261f2d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[15]));
  AL_DFF_X al_26a87873 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[16]));
  AL_DFF_X al_4ba6c514 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[17]));
  AL_DFF_X al_8483ed1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[0]));
  AL_DFF_X al_3c14f403 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[18]));
  AL_DFF_X al_d2a3a3ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[19]));
  AL_DFF_X al_2ee07a38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[20]));
  AL_DFF_X al_70c45082 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[21]));
  AL_DFF_X al_449f17bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[22]));
  AL_DFF_X al_dc01bb53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[23]));
  AL_DFF_X al_6dd2a1d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[24]));
  AL_DFF_X al_6de25d4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[25]));
  AL_DFF_X al_6b39c149 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[26]));
  AL_DFF_X al_a2ebe9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[27]));
  AL_DFF_X al_81452488 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[1]));
  AL_DFF_X al_6732ef46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[28]));
  AL_DFF_X al_89cf0a1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[29]));
  AL_DFF_X al_dea01056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[30]));
  AL_DFF_X al_3726bb4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[31]));
  AL_DFF_X al_e490898a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[2]));
  AL_DFF_X al_8e73cdf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[3]));
  AL_DFF_X al_753a51cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[4]));
  AL_DFF_X al_4bf2dbc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[5]));
  AL_DFF_X al_28bd37b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[6]));
  AL_DFF_X al_33df54b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6fd79ca[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fd032af[7]));
  AL_DFF_X al_97f2ae8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[8]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[8]));
  AL_DFF_X al_af8b35fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[9]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[9]));
  AL_DFF_X al_17598258 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[10]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[10]));
  AL_DFF_X al_c4382f68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[11]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[11]));
  AL_DFF_X al_236ad162 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[12]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[12]));
  AL_DFF_X al_9b44253 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[13]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[13]));
  AL_DFF_X al_4f556ebd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[14]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[14]));
  AL_DFF_X al_e26891db (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[15]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[15]));
  AL_DFF_X al_5175d6a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[16]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[16]));
  AL_DFF_X al_25943d39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[17]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[17]));
  AL_DFF_X al_5d993370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[18]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[18]));
  AL_DFF_X al_c6870073 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[19]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[19]));
  AL_DFF_X al_f2143f5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[20]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[20]));
  AL_DFF_X al_c81eb48c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[21]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[21]));
  AL_DFF_X al_948b4d8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[22]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[22]));
  AL_DFF_X al_d36e13c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[23]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[23]));
  AL_DFF_X al_c6a30bbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[24]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[24]));
  AL_DFF_X al_306b1c37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[25]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[25]));
  AL_DFF_X al_9e996eb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[26]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[26]));
  AL_DFF_X al_90c0a52b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[27]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[27]));
  AL_DFF_X al_3cdfcd24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[28]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[28]));
  AL_DFF_X al_40bcfc4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[29]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[29]));
  AL_DFF_X al_d8a36741 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[30]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[30]));
  AL_DFF_X al_7942aa3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[31]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[31]));
  AL_DFF_X al_1feccf0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[2]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[2]));
  AL_DFF_X al_4f6f2d05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[3]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[3]));
  AL_DFF_X al_56850569 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[4]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[4]));
  AL_DFF_X al_9d3458c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[5]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[5]));
  AL_DFF_X al_4151ad8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[6]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[6]));
  AL_DFF_X al_8de510b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[7]),
    .en(al_766b3b75),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c9327d6[7]));
  AL_DFF_X al_4e849cf9 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[8]));
  AL_DFF_X al_e99570e3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[9]));
  AL_DFF_X al_94baceb1 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[10]));
  AL_DFF_X al_a7bdadef (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[11]));
  AL_DFF_X al_8e59b7a3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[12]));
  AL_DFF_X al_82bb7642 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[13]));
  AL_DFF_X al_cf8c9b81 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[14]));
  AL_DFF_X al_61bc367d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[15]));
  AL_DFF_X al_7ddb34d8 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[16]));
  AL_DFF_X al_6fd277a9 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[17]));
  AL_DFF_X al_346cb299 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_271667bb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[0]));
  AL_DFF_X al_27549db7 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[18]));
  AL_DFF_X al_21ed2b79 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[19]));
  AL_DFF_X al_4a85e7e6 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[20]));
  AL_DFF_X al_7351c5f5 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[21]));
  AL_DFF_X al_20e8169 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[22]));
  AL_DFF_X al_d1f65a70 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[23]));
  AL_DFF_X al_6f45a97 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[24]));
  AL_DFF_X al_b27408d6 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[25]));
  AL_DFF_X al_1ec1b404 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[26]));
  AL_DFF_X al_83edb014 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[27]));
  AL_DFF_X al_386d10d2 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[1]));
  AL_DFF_X al_435e87d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[28]));
  AL_DFF_X al_9389602b (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[29]));
  AL_DFF_X al_1383530f (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[30]));
  AL_DFF_X al_e0e7f77a (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(al_bde0dc95[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[31]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(((E*C)*~(F)*~(B)+(E*C)*F*~(B)+~((E*C))*F*B+(E*C)*F*B))*~(A)+D*((E*C)*~(F)*~(B)+(E*C)*F*~(B)+~((E*C))*F*B+(E*C)*F*B)*~(A)+~(D)*((E*C)*~(F)*~(B)+(E*C)*F*~(B)+~((E*C))*F*B+(E*C)*F*B)*A+D*((E*C)*~(F)*~(B)+(E*C)*F*~(B)+~((E*C))*F*B+(E*C)*F*B)*A)"),
    .INIT(64'hfda8dd8875205500))
    al_3393c92b (
    .a(al_6f809586),
    .b(al_ee66e790),
    .c(al_53cc722d),
    .d(al_a16ef20a[0]),
    .e(al_ccabc055[0]),
    .f(al_4d016a39),
    .o(al_271667bb));
  AL_DFF_X al_83cae527 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[2]));
  AL_DFF_X al_910cd663 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[3]));
  AL_DFF_X al_94265a4 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[4]));
  AL_DFF_X al_bcfc8513 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[5]));
  AL_DFF_X al_68ceb98c (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[6]));
  AL_DFF_X al_f853697d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bde0dc95[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a16ef20a[7]));
  AL_DFF_X al_d7fc5dde (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[24]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[8]));
  AL_DFF_X al_4fbd101 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[25]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[9]));
  AL_DFF_X al_77b1fb98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[26]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[10]));
  AL_DFF_X al_8a9e7f14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[27]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[11]));
  AL_DFF_X al_f1614eef (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[28]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[12]));
  AL_DFF_X al_cc885919 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[29]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[13]));
  AL_DFF_X al_78bf20b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[30]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[14]));
  AL_DFF_X al_638f2cf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[31]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[15]));
  AL_DFF_X al_3103b6e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[16]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[0]));
  AL_DFF_X al_c9ca393 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[17]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[1]));
  AL_DFF_X al_be1f0c8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[18]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[2]));
  AL_DFF_X al_6a22527f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[19]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[3]));
  AL_DFF_X al_fdeb8a96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[20]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[4]));
  AL_DFF_X al_cf8fdd16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[21]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[5]));
  AL_DFF_X al_5bc0e012 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[22]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[6]));
  AL_DFF_X al_58a913c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_cf18c1c6[23]),
    .en(al_1d3bfd2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd02584[7]));
  AL_DFF_X al_773f9c71 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[8]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[8]));
  AL_DFF_X al_a48bb419 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[9]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[9]));
  AL_DFF_X al_bdc36a94 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[10]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[10]));
  AL_DFF_X al_f6235205 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[11]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[11]));
  AL_DFF_X al_fbcd425d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[12]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[12]));
  AL_DFF_X al_5f6a5375 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[13]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[13]));
  AL_DFF_X al_f4456fec (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[14]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[14]));
  AL_DFF_X al_cae9fe02 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[15]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[15]));
  AL_DFF_X al_fddb0724 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[16]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[16]));
  AL_DFF_X al_19f7cb25 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[17]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[17]));
  AL_DFF_X al_e4d92c09 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[18]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[18]));
  AL_DFF_X al_70348335 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[19]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[19]));
  AL_DFF_X al_28da7c5e (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[20]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[20]));
  AL_DFF_X al_100d30b3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[21]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[21]));
  AL_DFF_X al_ea1ee75c (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[22]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[22]));
  AL_DFF_X al_a758dcd2 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[23]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[23]));
  AL_DFF_X al_e14ede1f (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[24]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[24]));
  AL_DFF_X al_c1457613 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[25]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[25]));
  AL_DFF_X al_5f01547a (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[26]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[26]));
  AL_DFF_X al_6c56649e (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[27]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[27]));
  AL_DFF_X al_ecaca92d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[1]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[1]));
  AL_DFF_X al_1744ae49 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[28]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[28]));
  AL_DFF_X al_c175c62d (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[29]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[29]));
  AL_DFF_X al_d30fb1eb (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[30]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[30]));
  AL_DFF_X al_8c56da8f (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(al_c1211126[31]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[31]));
  AL_DFF_X al_212b2669 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[2]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[2]));
  AL_DFF_X al_dd82b6c1 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[3]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[3]));
  AL_DFF_X al_979c2af5 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[4]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[4]));
  AL_DFF_X al_f6868359 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[5]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[5]));
  AL_DFF_X al_e21f6722 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[6]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[6]));
  AL_DFF_X al_79fb3850 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c1211126[7]),
    .en(al_3f2c3141),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_126b3afd[7]));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~D*~(E*C*A)))"),
    .INIT(32'h33203300))
    al_97952e6b (
    .a(al_a8151162),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_c85db05d),
    .e(al_7b80e496[3]),
    .o(al_2dc65bff));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*C*A))"),
    .INIT(16'heccc))
    al_eba3db7f (
    .a(al_a8151162),
    .b(al_6ec8afa5),
    .c(al_a5849610),
    .d(al_7b80e496[2]),
    .o(al_2c78771b));
  AL_DFF_X al_e9db0f46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9d1d880c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b80e496[0]));
  AL_DFF_X al_6699da45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9d1d880c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b80e496[1]));
  AL_DFF_X al_9fbedd3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2c78771b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b80e496[2]));
  AL_DFF_X al_79b3f116 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2dc65bff),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7b80e496[3]));
  AL_DFF_X al_b08ad2a1 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c3eb1e82[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9b5530fd[0]));
  AL_DFF_X al_c186c1e0 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c3eb1e82[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9b5530fd[1]));
  AL_DFF_X al_64a545cd (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c3eb1e82[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9b5530fd[2]));
  AL_DFF_X al_76e218ab (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b537d840[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_202f2c67[0]));
  AL_DFF_X al_1cc15d04 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b537d840[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_202f2c67[1]));
  AL_DFF_X al_e5e8a3cc (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b537d840[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_202f2c67[2]));
  AL_DFF_X al_aadd51bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[8]));
  AL_DFF_X al_ff137e73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[9]));
  AL_DFF_X al_2bf9e3a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[10]));
  AL_DFF_X al_ec1e7eb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[11]));
  AL_DFF_X al_20a8629e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[12]));
  AL_DFF_X al_1293e58d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[13]));
  AL_DFF_X al_b7ba35d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[14]));
  AL_DFF_X al_28670d06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[15]));
  AL_DFF_X al_5c003cda (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[16]));
  AL_DFF_X al_aaa6a0cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[17]));
  AL_DFF_X al_1d927ed0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[0]));
  AL_DFF_X al_60ecf8da (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[18]));
  AL_DFF_X al_b17c748 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[19]));
  AL_DFF_X al_5aba3f95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[20]));
  AL_DFF_X al_8c6e2b2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[21]));
  AL_DFF_X al_b67c79a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[22]));
  AL_DFF_X al_20547503 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[23]));
  AL_DFF_X al_dc7b877f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[24]));
  AL_DFF_X al_1df2d7b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[25]));
  AL_DFF_X al_f14c4058 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[26]));
  AL_DFF_X al_1a16e7c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[27]));
  AL_DFF_X al_9414dc97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[1]));
  AL_DFF_X al_10f485e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[28]));
  AL_DFF_X al_71ec8417 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[29]));
  AL_DFF_X al_156ef330 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[30]));
  AL_DFF_X al_f868c0f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[31]));
  AL_DFF_X al_713c2d1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[2]));
  AL_DFF_X al_e3278660 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[3]));
  AL_DFF_X al_181c67ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[4]));
  AL_DFF_X al_26f28579 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[5]));
  AL_DFF_X al_34177cea (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[6]));
  AL_DFF_X al_924a611a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_1f3eaa15[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85a2bdb0[7]));
  AL_DFF_X al_af7e3546 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[8]));
  AL_DFF_X al_121c735b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[9]));
  AL_DFF_X al_f965d67f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[10]));
  AL_DFF_X al_77c6296a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[11]));
  AL_DFF_X al_6ba6a4a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[12]));
  AL_DFF_X al_88841dcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[13]));
  AL_DFF_X al_c0de9fdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[14]));
  AL_DFF_X al_878ef04a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[15]));
  AL_DFF_X al_3040536 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[16]));
  AL_DFF_X al_bcbe88e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[17]));
  AL_DFF_X al_38cdfba0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[0]));
  AL_DFF_X al_ff753ee6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[18]));
  AL_DFF_X al_d36a13dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[19]));
  AL_DFF_X al_8127a570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[20]));
  AL_DFF_X al_684b01b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[21]));
  AL_DFF_X al_ac2ec43a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[22]));
  AL_DFF_X al_baf3c5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[23]));
  AL_DFF_X al_a939715e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[24]));
  AL_DFF_X al_1a660ca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[25]));
  AL_DFF_X al_492aada2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[26]));
  AL_DFF_X al_53620619 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[27]));
  AL_DFF_X al_27e972f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[1]));
  AL_DFF_X al_7f07ea69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[28]));
  AL_DFF_X al_77d529e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[29]));
  AL_DFF_X al_68bd5cab (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[30]));
  AL_DFF_X al_6918d64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[31]));
  AL_DFF_X al_c0583a98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[2]));
  AL_DFF_X al_42b532b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[3]));
  AL_DFF_X al_495d4a20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[4]));
  AL_DFF_X al_935f1d3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[5]));
  AL_DFF_X al_2307a804 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[6]));
  AL_DFF_X al_ccc59fbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c7f68e2[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81a1940d[7]));
  AL_DFF_X al_8c0d10ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[8]));
  AL_DFF_X al_f7eb771c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[9]));
  AL_DFF_X al_94d8cfae (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[10]));
  AL_DFF_X al_54ef1332 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[11]));
  AL_DFF_X al_165875a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[12]));
  AL_DFF_X al_ee5cf9b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[13]));
  AL_DFF_X al_af75b7a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[14]));
  AL_DFF_X al_dcac7674 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[15]));
  AL_DFF_X al_42c2a940 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[16]));
  AL_DFF_X al_cf3fae4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[17]));
  AL_DFF_X al_cb83b621 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[0]));
  AL_DFF_X al_60b4401c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[18]));
  AL_DFF_X al_6e4325d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[19]));
  AL_DFF_X al_6bf98e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[20]));
  AL_DFF_X al_1353638a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[21]));
  AL_DFF_X al_7b99f32d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[22]));
  AL_DFF_X al_2d1da0cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[23]));
  AL_DFF_X al_c6ab3981 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[24]));
  AL_DFF_X al_fd1b3e52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[25]));
  AL_DFF_X al_93a1a61d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[26]));
  AL_DFF_X al_8a4f9feb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[27]));
  AL_DFF_X al_472998ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[1]));
  AL_DFF_X al_67dc47d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[28]));
  AL_DFF_X al_a72e3836 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[29]));
  AL_DFF_X al_6fb1aae8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[30]));
  AL_DFF_X al_3903b68a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[31]));
  AL_DFF_X al_a3f767f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[2]));
  AL_DFF_X al_7949e70f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[3]));
  AL_DFF_X al_7d01be47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[4]));
  AL_DFF_X al_fc11b7ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[5]));
  AL_DFF_X al_57f6b6d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[6]));
  AL_DFF_X al_2e3012dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8492e16[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe073fc9[7]));
  AL_DFF_X al_efdf58ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[8]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[8]));
  AL_DFF_X al_af14709e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[9]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[9]));
  AL_DFF_X al_bf075804 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[10]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[10]));
  AL_DFF_X al_ee42e75e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[11]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[11]));
  AL_DFF_X al_c4543f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[12]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[12]));
  AL_DFF_X al_c2c61477 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[13]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[13]));
  AL_DFF_X al_9a145c77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[14]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[14]));
  AL_DFF_X al_c0bc3b61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[15]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[15]));
  AL_DFF_X al_e7a96588 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[16]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[16]));
  AL_DFF_X al_fa95280b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[17]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[17]));
  AL_DFF_X al_3bbd9d48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f4b5275b),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[0]));
  AL_DFF_X al_43d686cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[18]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[18]));
  AL_DFF_X al_68a95d36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[19]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[19]));
  AL_DFF_X al_9b2b61d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[20]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[20]));
  AL_DFF_X al_703a0e34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[21]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[21]));
  AL_DFF_X al_b040a589 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[22]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[22]));
  AL_DFF_X al_c9a96958 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[23]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[23]));
  AL_DFF_X al_a8546243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[24]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[24]));
  AL_DFF_X al_57226817 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[25]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[25]));
  AL_DFF_X al_c7b1f011 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[26]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[26]));
  AL_DFF_X al_89190cbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[27]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[27]));
  AL_DFF_X al_9652e91c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2370214),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[1]));
  AL_DFF_X al_5ff8e1a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[28]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[28]));
  AL_DFF_X al_739c0744 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[29]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[29]));
  AL_DFF_X al_d6f71e72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[30]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[30]));
  AL_DFF_X al_2bde0dc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6e268dd3[31]),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[31]));
  AL_DFF_X al_432612ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bf952132),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[2]));
  AL_DFF_X al_bfe235ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_76a52f3d),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[3]));
  AL_DFF_X al_19b9c020 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c861c8f0),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[4]));
  AL_DFF_X al_38652411 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8a841cb4),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[5]));
  AL_DFF_X al_69595d30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_33a2911e),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[6]));
  AL_DFF_X al_f1fff8f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_73fb1ee5),
    .en(dBusAhb_HREADY_IN),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HWDATA[7]));
  AL_DFF_X al_582cabe4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_84a0e6),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bb6625de[0]));
  AL_DFF_X al_7fdbfd92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[12]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bb6625de[1]));
  AL_DFF_X al_c7154fcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c50e70c2),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1edb758f[0]));
  AL_DFF_X al_f7eaa42b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9ba628cf),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1edb758f[1]));
  AL_DFF_X al_bba93aff (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_40a6f08c[29]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_580ff8b7[0]));
  AL_DFF_X al_bd8f6d2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_40a6f08c[30]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_580ff8b7[1]));
  AL_MAP_LUT5 #(
    .EQN("(A*(C*B)*D*~(E)+~(A)*~((C*B))*~(D)*E+A*~((C*B))*~(D)*E+~(A)*(C*B)*~(D)*E+A*(C*B)*~(D)*E+A*~((C*B))*D*E+A*(C*B)*D*E)"),
    .INIT(32'haaff8000))
    al_ae872fde (
    .a(al_89ab45b5),
    .b(al_172eec6a),
    .c(al_a1a600b6),
    .d(al_ac1a4f11),
    .e(al_86d3f01a[2]),
    .o(al_25ff0fe3));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*(C*B)*D*~(E)+A*(C*B)*D*~(E)+~(A)*~((C*B))*~(D)*E+A*~((C*B))*~(D)*E+~(A)*(C*B)*~(D)*E+A*(C*B)*~(D)*E+A*~((C*B))*D*E+~(A)*(C*B)*D*E+A*(C*B)*D*E)"),
    .INIT(32'heaffc000))
    al_594685c6 (
    .a(al_4d82afcf),
    .b(al_da7f07ab),
    .c(al_8869249d),
    .d(al_ac1a4f11),
    .e(al_86d3f01a[3]),
    .o(al_d3323cee));
  AL_DFF_X al_970ec96b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25ff0fe3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86d3f01a[2]));
  AL_DFF_X al_3037f77f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d3323cee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86d3f01a[3]));
  AL_DFF_X al_1856317d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_eb46e9d2),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5f1afb5[0]));
  AL_DFF_X al_9959112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_40a6f08c[27]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5f1afb5[1]));
  AL_DFF_X al_7526da65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[8]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[8]));
  AL_DFF_X al_37ec4f8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[9]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[9]));
  AL_DFF_X al_8eb6b791 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[10]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[10]));
  AL_DFF_X al_27b82fbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[11]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[11]));
  AL_DFF_X al_1eec7b76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[13]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(dBusAhb_HSIZE[1]));
  AL_DFF_X al_57517970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[14]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[14]));
  AL_DFF_X al_3c59b07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[15]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[15]));
  AL_DFF_X al_e4728e11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[16]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[16]));
  AL_DFF_X al_fbe19c44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[17]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[17]));
  AL_DFF_X al_55b29daa (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[0]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[0]));
  AL_DFF_X al_10bd9edd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[18]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[18]));
  AL_DFF_X al_80e4fba0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[19]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[19]));
  AL_DFF_X al_1b03e023 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[20]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[20]));
  AL_DFF_X al_7b0c5096 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[21]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[21]));
  AL_DFF_X al_e30afaea (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[22]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[22]));
  AL_DFF_X al_37790c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[23]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[23]));
  AL_DFF_X al_c097b56b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[24]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[24]));
  AL_DFF_X al_f7129a92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[25]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[25]));
  AL_DFF_X al_40deb603 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[26]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[26]));
  AL_DFF_X al_5bd6b3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[27]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[27]));
  AL_DFF_X al_1d430310 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[1]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[1]));
  AL_DFF_X al_6d61b98c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[28]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[28]));
  AL_DFF_X al_1120e8f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[29]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[29]));
  AL_DFF_X al_250d018b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[30]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[30]));
  AL_DFF_X al_e151ed8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[31]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[31]));
  AL_DFF_X al_5f850675 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[2]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[2]));
  AL_DFF_X al_48ef55b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[3]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[3]));
  AL_DFF_X al_6f6ecdf2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[4]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[4]));
  AL_DFF_X al_b064b515 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[6]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[6]));
  AL_DFF_X al_1804d42f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_85a2bdb0[7]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e03b3126[7]));
  AL_DFF_X al_c0fa366b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[8]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[8]));
  AL_DFF_X al_a5451c97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[9]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[9]));
  AL_DFF_X al_4b72eeff (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[10]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[10]));
  AL_DFF_X al_48f93e18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[11]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[11]));
  AL_DFF_X al_522f26b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[12]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[12]));
  AL_DFF_X al_7bbe9177 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[13]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[13]));
  AL_DFF_X al_a2a8c215 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[14]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[14]));
  AL_DFF_X al_4a20c999 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[15]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[15]));
  AL_DFF_X al_d27779f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[16]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[16]));
  AL_DFF_X al_78e8fb31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[17]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[17]));
  AL_DFF_X al_50333221 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[0]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[0]));
  AL_DFF_X al_9058d3c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[18]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[18]));
  AL_DFF_X al_1aa49e07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[19]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[19]));
  AL_DFF_X al_ab4473cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[20]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[20]));
  AL_DFF_X al_9dde993d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[21]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[21]));
  AL_DFF_X al_bf7be43c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[22]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[22]));
  AL_DFF_X al_217b6ebc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[23]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[23]));
  AL_DFF_X al_56d2108f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[24]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[24]));
  AL_DFF_X al_53e533da (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[25]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[25]));
  AL_DFF_X al_11de2a0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[26]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[26]));
  AL_DFF_X al_684ed2e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[27]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[27]));
  AL_DFF_X al_d7245375 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[1]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[1]));
  AL_DFF_X al_8d823db (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[28]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[28]));
  AL_DFF_X al_9bbc681c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[29]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[29]));
  AL_DFF_X al_613bee42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[30]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[30]));
  AL_DFF_X al_aaa523c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[31]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[31]));
  AL_DFF_X al_36986146 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[2]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[2]));
  AL_DFF_X al_32a765a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[3]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[3]));
  AL_DFF_X al_8cc27260 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[4]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[4]));
  AL_DFF_X al_e27fa4a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[5]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[5]));
  AL_DFF_X al_204faf09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[6]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[6]));
  AL_DFF_X al_e8b50be7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a16ef20a[7]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9bf95cff[7]));
  AL_DFF_X al_173cc903 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[8]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[8]));
  AL_DFF_X al_b98fe8bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[9]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[9]));
  AL_DFF_X al_5823e9e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[10]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[10]));
  AL_DFF_X al_1a30e8b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[11]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[11]));
  AL_DFF_X al_2b35c232 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[12]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[12]));
  AL_DFF_X al_e3f63fda (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[13]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[13]));
  AL_DFF_X al_ca77fc3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[14]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[14]));
  AL_DFF_X al_1a6ec0ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[15]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[15]));
  AL_DFF_X al_5898c0cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[16]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[16]));
  AL_DFF_X al_2154775 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[17]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[17]));
  AL_DFF_X al_6fd283b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[0]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[0]));
  AL_DFF_X al_af1e3073 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[18]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[18]));
  AL_DFF_X al_d626f486 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[19]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[19]));
  AL_DFF_X al_2fc1a7fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[20]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[20]));
  AL_DFF_X al_2fd243b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[21]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[21]));
  AL_DFF_X al_6929cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[22]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[22]));
  AL_DFF_X al_bcd48a67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[23]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[23]));
  AL_DFF_X al_5ecc2c75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[24]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[24]));
  AL_DFF_X al_9dd0c48c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[25]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[25]));
  AL_DFF_X al_52347b8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[26]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[26]));
  AL_DFF_X al_ed086b8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[27]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[27]));
  AL_DFF_X al_d7cc8e41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[1]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[1]));
  AL_DFF_X al_c8ecce8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[28]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[28]));
  AL_DFF_X al_e7b16951 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[29]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[29]));
  AL_DFF_X al_a427052e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[30]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[30]));
  AL_DFF_X al_735b8603 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[31]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[31]));
  AL_DFF_X al_68392110 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[2]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[2]));
  AL_DFF_X al_f91db513 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[3]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[3]));
  AL_DFF_X al_ca3c0348 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[4]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[4]));
  AL_DFF_X al_4ca3743c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[5]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[5]));
  AL_DFF_X al_10191c31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[6]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[6]));
  AL_DFF_X al_65a95918 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bbc99cd7[7]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8074bdb[7]));
  AL_DFF_X al_d0dff042 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[8]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[8]));
  AL_DFF_X al_91808d7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[9]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[9]));
  AL_DFF_X al_4070afc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[10]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[10]));
  AL_DFF_X al_a572191f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[11]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[11]));
  AL_DFF_X al_9f57c998 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[12]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[12]));
  AL_DFF_X al_fa694b88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[13]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[13]));
  AL_DFF_X al_9695c37d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[14]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[14]));
  AL_DFF_X al_52af54d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[15]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[15]));
  AL_DFF_X al_cc808b7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[16]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[16]));
  AL_DFF_X al_4a1fcebd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[17]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[17]));
  AL_DFF_X al_df86e563 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[0]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[0]));
  AL_DFF_X al_a266b71e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[18]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[18]));
  AL_DFF_X al_81431268 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[19]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[19]));
  AL_DFF_X al_3857fa0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[20]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[20]));
  AL_DFF_X al_17352ffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[21]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[21]));
  AL_DFF_X al_4a07f3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[22]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[22]));
  AL_DFF_X al_1dfe4754 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[23]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[23]));
  AL_DFF_X al_477f727 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[24]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[24]));
  AL_DFF_X al_562af2e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[25]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[25]));
  AL_DFF_X al_57705321 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[26]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[26]));
  AL_DFF_X al_83986a28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[27]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[27]));
  AL_DFF_X al_df2f8fc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[1]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[1]));
  AL_DFF_X al_66b55c12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[28]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[28]));
  AL_DFF_X al_2a8035b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[29]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[29]));
  AL_DFF_X al_692eb5ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[30]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[30]));
  AL_DFF_X al_301f22e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[31]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[31]));
  AL_DFF_X al_6dccafc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[2]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[2]));
  AL_DFF_X al_5d45954f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[3]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[3]));
  AL_DFF_X al_65d9423e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[4]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[4]));
  AL_DFF_X al_d2fefc4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[5]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[5]));
  AL_DFF_X al_d7c9816d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[6]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[6]));
  AL_DFF_X al_bdadc03c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_52ea52d7[7]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f7928e2[7]));
  AL_DFF_X al_e33bddbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_17dd8854),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_27c2eb8[0]));
  AL_DFF_X al_7c82af16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c6966291[20]),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_27c2eb8[1]));
  AL_DFF_X al_38add109 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_40dcfa8c),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_555b0990[0]));
  AL_DFF_X al_a10941aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_4ab1b7b3),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_555b0990[1]));
  AL_DFF_X al_2fdb24d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_de0f70d9),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1e88c0c[0]));
  AL_DFF_X al_b2db2982 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a8c60ee7),
    .en(al_5a744f0f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a1e88c0c[1]));
  AL_DFF_X al_fa662140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[8]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[8]));
  AL_DFF_X al_d881108d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[9]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[9]));
  AL_DFF_X al_9948b503 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[10]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[10]));
  AL_DFF_X al_91426546 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[11]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[11]));
  AL_DFF_X al_d0fa0bb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[12]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[12]));
  AL_DFF_X al_8feb38f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[13]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[13]));
  AL_DFF_X al_78c9bc77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[14]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[14]));
  AL_DFF_X al_9c65f79b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[15]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[15]));
  AL_DFF_X al_d1e4fbdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[16]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[16]));
  AL_DFF_X al_67644c83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[17]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[17]));
  AL_DFF_X al_7f83533f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[18]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[18]));
  AL_DFF_X al_12df0c63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[19]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[19]));
  AL_DFF_X al_a9f88199 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[20]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[20]));
  AL_DFF_X al_2efee8d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[21]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[21]));
  AL_DFF_X al_f20380e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[22]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[22]));
  AL_DFF_X al_8fe4172b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[23]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[23]));
  AL_DFF_X al_27b89f70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[24]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[24]));
  AL_DFF_X al_97adb643 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[25]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[25]));
  AL_DFF_X al_275c0341 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[26]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[26]));
  AL_DFF_X al_3d67f07c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[27]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[27]));
  AL_DFF_X al_6fbd69e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[1]));
  AL_DFF_X al_7304c348 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[28]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[28]));
  AL_DFF_X al_94378828 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[29]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[29]));
  AL_DFF_X al_26c43eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[30]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[30]));
  AL_DFF_X al_6d0984b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[31]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[31]));
  AL_DFF_X al_27465486 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[2]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[2]));
  AL_DFF_X al_6a45ef68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[3]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[3]));
  AL_DFF_X al_6a9b122d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[4]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[4]));
  AL_DFF_X al_e59c9388 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[5]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[5]));
  AL_DFF_X al_70a8067b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[6]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[6]));
  AL_DFF_X al_7e4a7297 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f2fa5dc[7]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_46ea2d9f[7]));
  AL_DFF_X al_fc65d394 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b5f1afb5[0]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53188262[0]));
  AL_DFF_X al_a75336f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_b5f1afb5[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53188262[1]));
  AL_DFF_X al_b7ba0792 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e03b3126[8]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[8]));
  AL_DFF_X al_eb5ab5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e03b3126[9]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[9]));
  AL_DFF_X al_d745186a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e03b3126[10]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[10]));
  AL_DFF_X al_d2e7b1df (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e03b3126[11]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[11]));
  AL_DFF_X al_1835b904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_bb6625de[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[12]));
  AL_DFF_X al_fb4dab6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HSIZE[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[13]));
  AL_DFF_X al_fc7f2c73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e03b3126[14]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[14]));
  AL_DFF_X al_71c7c51d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e03b3126[28]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[28]));
  AL_DFF_X al_f72d8936 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e03b3126[29]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[29]));
  AL_DFF_X al_f2d5917 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e03b3126[7]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a0e6869c[7]));
  AL_DFF_X al_7ebcc32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HADDR[0]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50f87e49[0]));
  AL_DFF_X al_5c66e961 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(dBusAhb_HADDR[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50f87e49[1]));
  AL_DFF_X al_4d3c6ad9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[8]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[8]));
  AL_DFF_X al_aa082109 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[9]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[9]));
  AL_DFF_X al_f295ec37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[10]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[10]));
  AL_DFF_X al_1ec2056b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[11]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[11]));
  AL_DFF_X al_f205bc9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[12]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[12]));
  AL_DFF_X al_c66b13da (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[13]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[13]));
  AL_DFF_X al_b0f609a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[14]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[14]));
  AL_DFF_X al_5a958507 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[15]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[15]));
  AL_DFF_X al_524a0083 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[16]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[16]));
  AL_DFF_X al_9f6cad3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[17]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[17]));
  AL_DFF_X al_c74a6c35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[0]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[0]));
  AL_DFF_X al_8bf57a2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[18]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[18]));
  AL_DFF_X al_d255810a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[19]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[19]));
  AL_DFF_X al_9cc767c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[20]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[20]));
  AL_DFF_X al_90df0992 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[21]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[21]));
  AL_DFF_X al_3e3f6963 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[22]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[22]));
  AL_DFF_X al_c75c2dfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[23]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[23]));
  AL_DFF_X al_de329040 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[24]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[24]));
  AL_DFF_X al_937febe8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[25]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[25]));
  AL_DFF_X al_b4dde6e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[26]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[26]));
  AL_DFF_X al_e8cd59bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[27]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[27]));
  AL_DFF_X al_882f5706 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[1]));
  AL_DFF_X al_d7d8c4dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[28]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[28]));
  AL_DFF_X al_2e601caa (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[29]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[29]));
  AL_DFF_X al_22bfe3f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[30]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[30]));
  AL_DFF_X al_7c75801 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[31]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[31]));
  AL_DFF_X al_9595af9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[2]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[2]));
  AL_DFF_X al_6acc8b72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[3]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[3]));
  AL_DFF_X al_f1507e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[4]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[4]));
  AL_DFF_X al_5b34a992 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[5]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[5]));
  AL_DFF_X al_1987b65d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[6]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[6]));
  AL_DFF_X al_a69f0736 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9bf95cff[7]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e7cde15[7]));
  AL_DFF_X al_f2beca1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[8]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[8]));
  AL_DFF_X al_b450971a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[9]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[9]));
  AL_DFF_X al_244d384 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[10]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[10]));
  AL_DFF_X al_4108d82d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[11]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[11]));
  AL_DFF_X al_2ac5919 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[12]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[12]));
  AL_DFF_X al_124ab088 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[13]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[13]));
  AL_DFF_X al_67894bab (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[14]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[14]));
  AL_DFF_X al_61a661b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[15]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[15]));
  AL_DFF_X al_129005b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[16]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[16]));
  AL_DFF_X al_f8c7aecb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[17]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[17]));
  AL_DFF_X al_11a1b1a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[0]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[0]));
  AL_DFF_X al_872d5c3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[18]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[18]));
  AL_DFF_X al_2573cd87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[19]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[19]));
  AL_DFF_X al_42e94c34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[20]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[20]));
  AL_DFF_X al_9609356c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[21]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[21]));
  AL_DFF_X al_d3c0d18d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[22]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[22]));
  AL_DFF_X al_e01e365b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[23]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[23]));
  AL_DFF_X al_a3b107e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[24]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[24]));
  AL_DFF_X al_474e158a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[25]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[25]));
  AL_DFF_X al_9617f161 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[26]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[26]));
  AL_DFF_X al_bb010f86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[27]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[27]));
  AL_DFF_X al_17272ba5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[1]));
  AL_DFF_X al_de58e00f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[28]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[28]));
  AL_DFF_X al_1c184fa8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[29]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[29]));
  AL_DFF_X al_f8de40c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[30]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[30]));
  AL_DFF_X al_ed09f28d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[31]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[31]));
  AL_DFF_X al_f880a83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[2]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[2]));
  AL_DFF_X al_abed7f43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[3]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[3]));
  AL_DFF_X al_640aa117 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[4]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[4]));
  AL_DFF_X al_444f3914 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[5]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[5]));
  AL_DFF_X al_d689dd23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[6]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[6]));
  AL_DFF_X al_89f6ab54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8221e5ce[7]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfc96350[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .INIT(16'hf3e2))
    al_23e6abb0 (
    .a(al_bec39e4d),
    .b(al_5e275e81),
    .c(al_7b80e496[1]),
    .d(al_1a8c7c22[1]),
    .o(al_c2ce02d3));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .INIT(16'hf3e2))
    al_526d1aee (
    .a(al_bec39e4d),
    .b(al_5e275e81),
    .c(al_7b80e496[0]),
    .d(al_1a8c7c22[0]),
    .o(al_6be7ae97));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_2d122c09 (
    .a(al_bec39e4d),
    .b(al_5e275e81),
    .c(al_7b80e496[2]),
    .d(al_86d3f01a[2]),
    .e(al_1a8c7c22[2]),
    .o(al_fdcd8a4d));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_7acbe7f3 (
    .a(al_bec39e4d),
    .b(al_5e275e81),
    .c(al_7b80e496[3]),
    .d(al_86d3f01a[3]),
    .e(al_1a8c7c22[3]),
    .o(al_92a03ec7));
  AL_DFF_X al_26f239a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6be7ae97),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1a8c7c22[0]));
  AL_DFF_X al_d9ef719d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c2ce02d3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1a8c7c22[1]));
  AL_DFF_X al_19f72465 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_fdcd8a4d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1a8c7c22[2]));
  AL_DFF_X al_5ff83783 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_92a03ec7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1a8c7c22[3]));
  AL_DFF_X al_7789eb6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_27c2eb8[0]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_727d2e98[0]));
  AL_DFF_X al_3f37be2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_27c2eb8[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_727d2e98[1]));
  AL_DFF_X al_391e2d37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[8]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[8]));
  AL_DFF_X al_30e905c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[9]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[9]));
  AL_DFF_X al_6389391f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[10]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[10]));
  AL_DFF_X al_b1ae6862 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[11]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[11]));
  AL_DFF_X al_957f9ce5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[12]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[12]));
  AL_DFF_X al_3938f4ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[13]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[13]));
  AL_DFF_X al_742a6834 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[14]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[14]));
  AL_DFF_X al_f7def0c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[15]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[15]));
  AL_DFF_X al_6a60d755 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[16]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[16]));
  AL_DFF_X al_fa1865f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[17]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[17]));
  AL_DFF_X al_aa6477a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[0]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[0]));
  AL_DFF_X al_e99b4a51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[18]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[18]));
  AL_DFF_X al_750bfd1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[19]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[19]));
  AL_DFF_X al_199415ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[20]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[20]));
  AL_DFF_X al_dd110adc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[21]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[21]));
  AL_DFF_X al_9a5eb3b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[22]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[22]));
  AL_DFF_X al_85e54ead (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[23]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[23]));
  AL_DFF_X al_91010185 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[24]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[24]));
  AL_DFF_X al_5a9e58ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[25]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[25]));
  AL_DFF_X al_43b10dae (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[26]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[26]));
  AL_DFF_X al_652696cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[27]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[27]));
  AL_DFF_X al_af523ac2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[1]));
  AL_DFF_X al_f4f68452 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[28]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[28]));
  AL_DFF_X al_d8746d2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[29]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[29]));
  AL_DFF_X al_461b4794 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[30]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[30]));
  AL_DFF_X al_5bf9b8ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[31]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[31]));
  AL_DFF_X al_1c01345e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[2]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[2]));
  AL_DFF_X al_34350c3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[3]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[3]));
  AL_DFF_X al_7a1b987a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[4]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[4]));
  AL_DFF_X al_92867dca (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[5]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[5]));
  AL_DFF_X al_2f200ffc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[6]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[6]));
  AL_DFF_X al_6cc19ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_9e82589f[7]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1fb6e0a[7]));
  AL_DFF_X al_cff1e2d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[8]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[8]));
  AL_DFF_X al_a2e7fc29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[9]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[9]));
  AL_DFF_X al_dce34a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[10]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[10]));
  AL_DFF_X al_7e4285ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[11]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[11]));
  AL_DFF_X al_1d95a0c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[12]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[12]));
  AL_DFF_X al_6bd1ef6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[13]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[13]));
  AL_DFF_X al_180a2599 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[14]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[14]));
  AL_DFF_X al_dcfcc450 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[15]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[15]));
  AL_DFF_X al_cd4afcff (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[16]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[16]));
  AL_DFF_X al_9c76eb1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[17]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[17]));
  AL_DFF_X al_8f08cb9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[0]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[0]));
  AL_DFF_X al_47a2d5d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[18]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[18]));
  AL_DFF_X al_491e8a09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[19]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[19]));
  AL_DFF_X al_7fcffb8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[20]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[20]));
  AL_DFF_X al_d676ea3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[21]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[21]));
  AL_DFF_X al_33f4bad3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[22]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[22]));
  AL_DFF_X al_14047f31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[23]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[23]));
  AL_DFF_X al_3c22a61c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[24]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[24]));
  AL_DFF_X al_b1e6690c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[25]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[25]));
  AL_DFF_X al_aa412121 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[26]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[26]));
  AL_DFF_X al_2afbe7ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[27]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[27]));
  AL_DFF_X al_42532176 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[1]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[1]));
  AL_DFF_X al_fcf74f05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[28]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[28]));
  AL_DFF_X al_dd213dac (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[29]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[29]));
  AL_DFF_X al_519602e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[30]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[30]));
  AL_DFF_X al_f069f098 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[31]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[31]));
  AL_DFF_X al_24c75df7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[2]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[2]));
  AL_DFF_X al_ef1dc479 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[3]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[3]));
  AL_DFF_X al_20a67f25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[4]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[4]));
  AL_DFF_X al_17d16b93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[5]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[5]));
  AL_DFF_X al_a099f3e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[6]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[6]));
  AL_DFF_X al_127027c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_830b3656[7]),
    .en(al_a430e4d2),
    .sr(~al_98842338),
    .ss(1'b0),
    .q(al_7b59c46e[7]));
  AL_DFF_X al_61a0fa03 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2d4f70b0[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d392f4f[0]));
  AL_DFF_X al_f8ff3336 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2d4f70b0[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d392f4f[1]));
  AL_DFF_X al_bcc82701 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2d4f70b0[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d392f4f[2]));
  AL_DFF_X al_30b8896a (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2d4f70b0[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d392f4f[3]));
  AL_DFF_X al_333b6655 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2d4f70b0[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d392f4f[4]));
  AL_DFF_X al_155d2111 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2d4f70b0[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d392f4f[5]));
  AL_DFF_X al_9db3d031 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[8]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[8]));
  AL_DFF_X al_51b4fa4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[9]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[9]));
  AL_DFF_X al_f42c4388 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[10]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[10]));
  AL_DFF_X al_3dbc12db (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[11]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[11]));
  AL_DFF_X al_fb8e96c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[12]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[12]));
  AL_DFF_X al_cc5c71b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[13]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[13]));
  AL_DFF_X al_81297cae (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[14]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[14]));
  AL_DFF_X al_bb8b3df5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[15]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[15]));
  AL_DFF_X al_17e9d5f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[16]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[16]));
  AL_DFF_X al_a73353bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[17]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[17]));
  AL_DFF_X al_bf515542 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_94f1da4c[0]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[0]));
  AL_DFF_X al_4555bad1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[18]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[18]));
  AL_DFF_X al_b4fee469 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[19]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[19]));
  AL_DFF_X al_7ae81728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[20]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[20]));
  AL_DFF_X al_5d02d63e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[21]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[21]));
  AL_DFF_X al_18897cc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[22]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[22]));
  AL_DFF_X al_88931c76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[23]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[23]));
  AL_DFF_X al_4094be5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[24]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[24]));
  AL_DFF_X al_74569fa5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[25]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[25]));
  AL_DFF_X al_938c1a70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[26]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[26]));
  AL_DFF_X al_2257dfdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[27]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[27]));
  AL_DFF_X al_d173e0ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[1]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[1]));
  AL_DFF_X al_56825126 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[28]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[28]));
  AL_DFF_X al_af940374 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[29]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[29]));
  AL_DFF_X al_20ea28e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[30]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[30]));
  AL_DFF_X al_c0081590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[31]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[31]));
  AL_DFF_X al_70a7a49c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[2]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[2]));
  AL_DFF_X al_6e08612b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[3]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[3]));
  AL_DFF_X al_73e6e1ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[4]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[4]));
  AL_DFF_X al_4c354f41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[5]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[5]));
  AL_DFF_X al_1c753898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[6]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[6]));
  AL_DFF_X al_19d64476 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_32172a12[7]),
    .en(al_3f04848f),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec26021c[7]));
  AL_DFF_X al_a6559e2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[8]));
  AL_DFF_X al_7bfaae22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[9]));
  AL_DFF_X al_6e646313 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[10]));
  AL_DFF_X al_f7cd7493 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[11]));
  AL_DFF_X al_95a78603 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[12]));
  AL_DFF_X al_885e7594 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[13]));
  AL_DFF_X al_d9920508 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[14]));
  AL_DFF_X al_c3374a25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[15]));
  AL_DFF_X al_a5e9e08a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[16]));
  AL_DFF_X al_519ee93c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[17]));
  AL_DFF_X al_53be9e02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[0]));
  AL_DFF_X al_1ff6ab6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[18]));
  AL_DFF_X al_90f30d03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[19]));
  AL_DFF_X al_2906140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[20]));
  AL_DFF_X al_94814473 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[21]));
  AL_DFF_X al_d8bfa0a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[22]));
  AL_DFF_X al_913530d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[23]));
  AL_DFF_X al_df300068 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[24]));
  AL_DFF_X al_de617911 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[25]));
  AL_DFF_X al_e446dcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[26]));
  AL_DFF_X al_92261327 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[27]));
  AL_DFF_X al_8ee55a7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[1]));
  AL_DFF_X al_3767b345 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[28]));
  AL_DFF_X al_903dae36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[29]));
  AL_DFF_X al_3ca5d926 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[30]));
  AL_DFF_X al_77de8e16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[31]));
  AL_DFF_X al_94207e8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[2]));
  AL_DFF_X al_e4caec90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[3]));
  AL_DFF_X al_1e201e1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[4]));
  AL_DFF_X al_25e37a50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[5]));
  AL_DFF_X al_dcc548a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[6]));
  AL_DFF_X al_1d929d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_d0c02c51[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b70cb9be[7]));
  AL_DFF_X al_4eb041e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[8]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[8]));
  AL_DFF_X al_ba96267 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[9]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[9]));
  AL_DFF_X al_cf0d7128 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[10]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[10]));
  AL_DFF_X al_d1381672 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[11]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[11]));
  AL_DFF_X al_99bc4f07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[12]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[12]));
  AL_DFF_X al_1242dc24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[13]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[13]));
  AL_DFF_X al_f3bacbaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[14]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[14]));
  AL_DFF_X al_5704823 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[15]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[15]));
  AL_DFF_X al_338964a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[16]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[16]));
  AL_DFF_X al_6fb20cae (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[17]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[17]));
  AL_DFF_X al_4641986c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f4b5275b),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[0]));
  AL_DFF_X al_e4ffb375 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[18]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[18]));
  AL_DFF_X al_d6a291a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[19]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[19]));
  AL_DFF_X al_c5c3b52f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[20]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[20]));
  AL_DFF_X al_e5364bf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[21]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[21]));
  AL_DFF_X al_aa7b09c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[22]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[22]));
  AL_DFF_X al_53f32607 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[23]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[23]));
  AL_DFF_X al_43310da3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[24]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[24]));
  AL_DFF_X al_664afb6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[25]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[25]));
  AL_DFF_X al_2384fac1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[26]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[26]));
  AL_DFF_X al_4479aed (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[27]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[27]));
  AL_DFF_X al_935be2b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[1]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[1]));
  AL_DFF_X al_9a032585 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[28]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[28]));
  AL_DFF_X al_ffc230fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[29]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[29]));
  AL_DFF_X al_a43ba6eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[30]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[30]));
  AL_DFF_X al_82740ccb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[31]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[31]));
  AL_DFF_X al_6857e0d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[2]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[2]));
  AL_DFF_X al_d2d0da34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[3]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[3]));
  AL_DFF_X al_b3ebcbdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[4]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[4]));
  AL_DFF_X al_2ffa14d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[5]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[5]));
  AL_DFF_X al_2fac98c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[6]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[6]));
  AL_DFF_X al_323e02ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_f337bb3c[7]),
    .en(al_bb0cd305),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f12834e3[7]));
  AL_DFF_X al_7539b08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_53188262[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_212ac3ba[0]));
  AL_DFF_X al_42a4d67f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_53188262[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_212ac3ba[1]));
  AL_DFF_X al_e6b277a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[8]));
  AL_DFF_X al_d8127c6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[9]));
  AL_DFF_X al_52777016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[10]));
  AL_DFF_X al_a3a39d6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[11]));
  AL_DFF_X al_c74e4b9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[12]));
  AL_DFF_X al_b27c2d73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[13]));
  AL_DFF_X al_db2b0e71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[14]));
  AL_DFF_X al_e1d41f02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[28]));
  AL_DFF_X al_11835682 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[29]));
  AL_DFF_X al_2e62d096 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a0e6869c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36a894af[7]));
  AL_DFF_X al_368c8f8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_50f87e49[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70c1ae82[0]));
  AL_DFF_X al_c2c73691 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_50f87e49[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70c1ae82[1]));
  AL_DFF_X al_df3fb297 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[8]));
  AL_DFF_X al_294995e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[9]));
  AL_DFF_X al_6f083f7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[10]));
  AL_DFF_X al_2b81b99f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[11]));
  AL_DFF_X al_92585a0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[12]));
  AL_DFF_X al_5a849634 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[13]));
  AL_DFF_X al_526080d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[14]));
  AL_DFF_X al_9fabf20b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[15]));
  AL_DFF_X al_e6d27cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[16]));
  AL_DFF_X al_58461eeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[17]));
  AL_DFF_X al_bd311eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[0]));
  AL_DFF_X al_351916f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[18]));
  AL_DFF_X al_c8384fda (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[19]));
  AL_DFF_X al_38112e64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[20]));
  AL_DFF_X al_73c5f3d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[21]));
  AL_DFF_X al_fc33920a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[22]));
  AL_DFF_X al_1baa7011 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[23]));
  AL_DFF_X al_e74ca2bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[24]));
  AL_DFF_X al_3a3efe4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[25]));
  AL_DFF_X al_70b90f5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[26]));
  AL_DFF_X al_2ea97875 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[27]));
  AL_DFF_X al_f67c728c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[1]));
  AL_DFF_X al_7f032f1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[28]));
  AL_DFF_X al_5a781b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[29]));
  AL_DFF_X al_5b24994b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[30]));
  AL_DFF_X al_b0d2b61b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_72cf1502),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[31]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_5a26d42a (
    .a(dBusAhb_HRDATA[31]),
    .b(al_aabf3e05),
    .o(al_72cf1502));
  AL_DFF_X al_b559c8be (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[2]));
  AL_DFF_X al_800c413d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[3]));
  AL_DFF_X al_56eb3ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[4]));
  AL_DFF_X al_406f4408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[5]));
  AL_DFF_X al_7b4968fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[6]));
  AL_DFF_X al_86bf6afb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8c4e5d9c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_24ce3017[7]));
  AL_DFF_X al_9a460b9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[8]));
  AL_DFF_X al_3cc714e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[9]));
  AL_DFF_X al_b3d79fbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[10]));
  AL_DFF_X al_e12f50be (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[11]));
  AL_DFF_X al_9c9db9a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[12]));
  AL_DFF_X al_f556966d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[13]));
  AL_DFF_X al_e38932af (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[14]));
  AL_DFF_X al_77b691cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[15]));
  AL_DFF_X al_ca703101 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[16]));
  AL_DFF_X al_27d0be38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[17]));
  AL_DFF_X al_329a8f86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[0]));
  AL_DFF_X al_c9f7cf57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[18]));
  AL_DFF_X al_54fa6da3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[19]));
  AL_DFF_X al_ec70afdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[20]));
  AL_DFF_X al_8d493aea (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[21]));
  AL_DFF_X al_ae803213 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[22]));
  AL_DFF_X al_ab943338 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[23]));
  AL_DFF_X al_e5295963 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[24]));
  AL_DFF_X al_209954fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[25]));
  AL_DFF_X al_31572404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[26]));
  AL_DFF_X al_61cc19a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[27]));
  AL_DFF_X al_162feea4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[1]));
  AL_DFF_X al_d4a91932 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[28]));
  AL_DFF_X al_6dada6c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[29]));
  AL_DFF_X al_db9e1d43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[30]));
  AL_DFF_X al_42c449ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[31]));
  AL_DFF_X al_a9dd1edd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[32]));
  AL_DFF_X al_90974a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[33]));
  AL_DFF_X al_534ee505 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[34]));
  AL_DFF_X al_8ad90af5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[35]));
  AL_DFF_X al_8a8e927e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[36]));
  AL_DFF_X al_416b5a4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[37]));
  AL_DFF_X al_9bb62b2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[2]));
  AL_DFF_X al_eaca7dd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[38]));
  AL_DFF_X al_77871d50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[39]));
  AL_DFF_X al_1dc84940 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[40]));
  AL_DFF_X al_5fb51be0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[41]));
  AL_DFF_X al_4144b9c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[42]));
  AL_DFF_X al_1a582d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[43]));
  AL_DFF_X al_4b4cd1bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[44]));
  AL_DFF_X al_77673509 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[45]));
  AL_DFF_X al_b530baa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[46]));
  AL_DFF_X al_528735d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[47]));
  AL_DFF_X al_96f67265 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[3]));
  AL_DFF_X al_72b753b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[48]));
  AL_DFF_X al_a753aa28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[49]));
  AL_DFF_X al_43ff2c31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[50]));
  AL_DFF_X al_94798b5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8dd2d746[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[51]));
  AL_DFF_X al_90887a81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[4]));
  AL_DFF_X al_cd302338 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[5]));
  AL_DFF_X al_7584caab (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[6]));
  AL_DFF_X al_a9ff7c97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_ccb50b3a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71c7f8f0[7]));
  AL_DFF_X al_cac20196 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[8]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[8]));
  AL_DFF_X al_6669ccb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[9]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[9]));
  AL_DFF_X al_1854dccf (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[10]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[10]));
  AL_DFF_X al_600f2f29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[11]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[11]));
  AL_DFF_X al_81785080 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[12]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[12]));
  AL_DFF_X al_db1b08a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[13]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[13]));
  AL_DFF_X al_7686afb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[14]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[14]));
  AL_DFF_X al_7dfc7cdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[15]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[15]));
  AL_DFF_X al_a8e7e842 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[16]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[16]));
  AL_DFF_X al_3959d1df (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[17]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[17]));
  AL_DFF_X al_5bcb81c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[0]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[0]));
  AL_DFF_X al_7ef47a57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[18]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[18]));
  AL_DFF_X al_c9132a26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[19]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[19]));
  AL_DFF_X al_84c12a0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[20]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[20]));
  AL_DFF_X al_f37c990d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[21]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[21]));
  AL_DFF_X al_160e1608 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[22]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[22]));
  AL_DFF_X al_bfebf86a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[23]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[23]));
  AL_DFF_X al_86cee06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[24]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[24]));
  AL_DFF_X al_7e2d4bc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[25]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[25]));
  AL_DFF_X al_5aed53fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[26]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[26]));
  AL_DFF_X al_7fea0d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[27]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[27]));
  AL_DFF_X al_b8673911 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[1]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[1]));
  AL_DFF_X al_c42bb4e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[28]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[28]));
  AL_DFF_X al_c931277a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[29]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[29]));
  AL_DFF_X al_3cc3512f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[30]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[30]));
  AL_DFF_X al_b0f2e7f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[31]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[31]));
  AL_DFF_X al_c2cc8b8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[2]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[2]));
  AL_DFF_X al_94597cfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[3]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[3]));
  AL_DFF_X al_c4496e54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[4]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[4]));
  AL_DFF_X al_c6ba05ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[5]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[5]));
  AL_DFF_X al_494d53ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[6]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[6]));
  AL_DFF_X al_4869887f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_2e7cde15[7]),
    .en(al_99763382),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e45b51d9[7]));
  AL_DFF_X al_c468b8d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[8]));
  AL_DFF_X al_89e26a77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[9]));
  AL_DFF_X al_868d72ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[10]));
  AL_DFF_X al_2a0c699d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[11]));
  AL_DFF_X al_747d0f52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[12]));
  AL_DFF_X al_bf0c5c3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[13]));
  AL_DFF_X al_96e630ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[14]));
  AL_DFF_X al_652545dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[15]));
  AL_DFF_X al_77370b43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[16]));
  AL_DFF_X al_84d9f4fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[17]));
  AL_DFF_X al_c0b83f20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[0]));
  AL_DFF_X al_1a50717 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[18]));
  AL_DFF_X al_ecaf1fe5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[19]));
  AL_DFF_X al_b8ab2c7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[20]));
  AL_DFF_X al_4be11b07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[21]));
  AL_DFF_X al_9f9bf732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[22]));
  AL_DFF_X al_b7de97e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[23]));
  AL_DFF_X al_3e17b913 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[24]));
  AL_DFF_X al_26921b5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[25]));
  AL_DFF_X al_f7bdb28c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[26]));
  AL_DFF_X al_5ff8787f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[27]));
  AL_DFF_X al_403b4c6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[1]));
  AL_DFF_X al_be4dac9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[28]));
  AL_DFF_X al_fd7831f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[29]));
  AL_DFF_X al_5eab5e25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[30]));
  AL_DFF_X al_48925f80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[31]));
  AL_DFF_X al_f9a3c587 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[2]));
  AL_DFF_X al_e075bae3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[3]));
  AL_DFF_X al_82374f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[4]));
  AL_DFF_X al_a60fa4e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[5]));
  AL_DFF_X al_5c95831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[6]));
  AL_DFF_X al_be3f5d17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8aeaa5c1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8900fb4e[7]));
  AL_DFF_X al_2d332181 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_74dc1091[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c72a609[0]));
  AL_DFF_X al_a161bd6e (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_74dc1091[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c72a609[1]));
  AL_DFF_X al_53d92684 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_74dc1091[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c72a609[2]));
  AL_DFF_X al_8a8b16d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[8]));
  AL_DFF_X al_d727f9b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[9]));
  AL_DFF_X al_7e3a21c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[10]));
  AL_DFF_X al_3760c928 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[11]));
  AL_DFF_X al_13002661 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[12]));
  AL_DFF_X al_897c57e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[13]));
  AL_DFF_X al_4022b915 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[14]));
  AL_DFF_X al_e7377164 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[15]));
  AL_DFF_X al_34e562cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[16]));
  AL_DFF_X al_fc467db6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[17]));
  AL_DFF_X al_33dac670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[0]));
  AL_DFF_X al_892ea019 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[18]));
  AL_DFF_X al_74ee1da3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[19]));
  AL_DFF_X al_a486f839 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[20]));
  AL_DFF_X al_808b89fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[21]));
  AL_DFF_X al_d9dce85c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[22]));
  AL_DFF_X al_dde1385f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[23]));
  AL_DFF_X al_54afac3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[24]));
  AL_DFF_X al_85c9e91f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[25]));
  AL_DFF_X al_ed846d8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[26]));
  AL_DFF_X al_412d2ae5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[27]));
  AL_DFF_X al_83b0a70a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[1]));
  AL_DFF_X al_34796d85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[28]));
  AL_DFF_X al_d2e9f2ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[29]));
  AL_DFF_X al_e269cdb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[30]));
  AL_DFF_X al_25eabbca (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[31]));
  AL_DFF_X al_63fc9b90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[2]));
  AL_DFF_X al_8dffbf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[3]));
  AL_DFF_X al_13268b96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[4]));
  AL_DFF_X al_14d3140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[5]));
  AL_DFF_X al_c54a97a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[6]));
  AL_DFF_X al_1f09422d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c28c3a52[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccabc055[7]));
  AL_DFF_X al_6c877aee (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(al_591b5570[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12792818[0]));
  AL_DFF_X al_f4fabf36 (
    .ar(1'b0),
    .as(SYS_RST_o),
    .clk(SYS_CLK),
    .d(al_591b5570[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12792818[1]));
  AL_DFF_X al_82d79944 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[8]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[8]));
  AL_DFF_X al_23db2e97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[9]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[9]));
  AL_DFF_X al_ad2b242d (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[10]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[10]));
  AL_DFF_X al_4f6f2b6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[11]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[11]));
  AL_DFF_X al_2d7cd930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[12]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[12]));
  AL_DFF_X al_c792e427 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[13]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[13]));
  AL_DFF_X al_37703eb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[14]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[14]));
  AL_DFF_X al_8b3e11ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[15]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[15]));
  AL_DFF_X al_694b073e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[16]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[16]));
  AL_DFF_X al_c0203ca2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[17]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[17]));
  AL_DFF_X al_9b0f7a05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[0]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[0]));
  AL_DFF_X al_e8877170 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[18]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[18]));
  AL_DFF_X al_d63a8bc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[19]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[19]));
  AL_DFF_X al_6f25cf47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[20]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[20]));
  AL_DFF_X al_55549ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[21]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[21]));
  AL_DFF_X al_f88d5744 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[22]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[22]));
  AL_DFF_X al_8f171db9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[23]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[23]));
  AL_DFF_X al_77a036ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[24]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[24]));
  AL_DFF_X al_16f4f2cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[25]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[25]));
  AL_DFF_X al_4e09062e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[26]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[26]));
  AL_DFF_X al_a05d34cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[27]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[27]));
  AL_DFF_X al_8b587c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[1]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[1]));
  AL_DFF_X al_aadb8779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[28]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[28]));
  AL_DFF_X al_bc938e21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[29]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[29]));
  AL_DFF_X al_5f2e7601 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[30]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[30]));
  AL_DFF_X al_cac73619 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[31]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[31]));
  AL_DFF_X al_77bcbfd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[2]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[2]));
  AL_DFF_X al_b33323fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[3]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[3]));
  AL_DFF_X al_9b56774 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[4]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[4]));
  AL_DFF_X al_239b78b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[5]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[5]));
  AL_DFF_X al_97dc0e8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[6]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[6]));
  AL_DFF_X al_a4677ead (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_45e5d9f7[7]),
    .en(al_5e275e81),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97943858[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_221c1845 (
    .a(1'b0),
    .o({al_22240f9f,open_n108}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e4508536 (
    .a(al_7b59c46e[7]),
    .b(al_f12834e3[8]),
    .c(al_91974942),
    .o({al_d135ca94,al_a5f7e6c[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8d01ba9d (
    .a(al_7b59c46e[8]),
    .b(al_f12834e3[9]),
    .c(al_d135ca94),
    .o({al_ab9e30a4,al_a5f7e6c[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9355ef8d (
    .a(al_7b59c46e[9]),
    .b(al_f12834e3[10]),
    .c(al_ab9e30a4),
    .o({al_4d279efb,al_a5f7e6c[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_73c453a5 (
    .a(al_7b59c46e[10]),
    .b(al_f12834e3[11]),
    .c(al_4d279efb),
    .o({al_ae1b5d59,al_a5f7e6c[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_acac78ae (
    .a(al_7b59c46e[11]),
    .b(al_f12834e3[12]),
    .c(al_ae1b5d59),
    .o({al_f466006e,al_a5f7e6c[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_76b50717 (
    .a(al_7b59c46e[12]),
    .b(al_f12834e3[13]),
    .c(al_f466006e),
    .o({al_4d64c75,al_a5f7e6c[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3f3743ea (
    .a(al_7b59c46e[13]),
    .b(al_f12834e3[14]),
    .c(al_4d64c75),
    .o({al_5a617f02,al_a5f7e6c[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_726182ce (
    .a(al_7b59c46e[14]),
    .b(al_f12834e3[15]),
    .c(al_5a617f02),
    .o({al_c63a3306,al_a5f7e6c[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eda24893 (
    .a(al_7b59c46e[15]),
    .b(al_f12834e3[16]),
    .c(al_c63a3306),
    .o({al_6b46d3b9,al_a5f7e6c[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_123b9aab (
    .a(al_7b59c46e[16]),
    .b(al_f12834e3[17]),
    .c(al_6b46d3b9),
    .o({al_8c8f6789,al_a5f7e6c[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2cd0a58e (
    .a(al_b70cb9be[31]),
    .b(al_f12834e3[0]),
    .c(al_22240f9f),
    .o({al_e9e54e67,al_a5f7e6c[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4e48b126 (
    .a(al_7b59c46e[17]),
    .b(al_f12834e3[18]),
    .c(al_8c8f6789),
    .o({al_443b56a1,al_a5f7e6c[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b76fdfa3 (
    .a(al_7b59c46e[18]),
    .b(al_f12834e3[19]),
    .c(al_443b56a1),
    .o({al_19286ed8,al_a5f7e6c[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b2492cd (
    .a(al_7b59c46e[19]),
    .b(al_f12834e3[20]),
    .c(al_19286ed8),
    .o({al_82a462e4,al_a5f7e6c[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2a170320 (
    .a(al_7b59c46e[20]),
    .b(al_f12834e3[21]),
    .c(al_82a462e4),
    .o({al_2f093a42,al_a5f7e6c[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b48f290a (
    .a(al_7b59c46e[21]),
    .b(al_f12834e3[22]),
    .c(al_2f093a42),
    .o({al_debb551a,al_a5f7e6c[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1a4c9947 (
    .a(al_7b59c46e[22]),
    .b(al_f12834e3[23]),
    .c(al_debb551a),
    .o({al_cd5a3103,al_a5f7e6c[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d786296 (
    .a(al_7b59c46e[23]),
    .b(al_f12834e3[24]),
    .c(al_cd5a3103),
    .o({al_24003c83,al_a5f7e6c[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f0b5c006 (
    .a(al_7b59c46e[24]),
    .b(al_f12834e3[25]),
    .c(al_24003c83),
    .o({al_ec08a0e6,al_a5f7e6c[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_18a8f8a7 (
    .a(al_7b59c46e[25]),
    .b(al_f12834e3[26]),
    .c(al_ec08a0e6),
    .o({al_c06b4d62,al_a5f7e6c[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_42f32459 (
    .a(al_7b59c46e[26]),
    .b(al_f12834e3[27]),
    .c(al_c06b4d62),
    .o({al_c862b555,al_a5f7e6c[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_37c675ff (
    .a(al_7b59c46e[0]),
    .b(al_f12834e3[1]),
    .c(al_e9e54e67),
    .o({al_dfe2f2a3,al_a5f7e6c[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d941e571 (
    .a(al_7b59c46e[27]),
    .b(al_f12834e3[28]),
    .c(al_c862b555),
    .o({al_c28f9c66,al_a5f7e6c[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b743a90 (
    .a(al_7b59c46e[28]),
    .b(al_f12834e3[29]),
    .c(al_c28f9c66),
    .o({al_3f573e25,al_a5f7e6c[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_25a7fcce (
    .a(al_7b59c46e[29]),
    .b(al_f12834e3[30]),
    .c(al_3f573e25),
    .o({al_62997e0b,al_a5f7e6c[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6b49ebdb (
    .a(al_7b59c46e[30]),
    .b(al_f12834e3[31]),
    .c(al_62997e0b),
    .o({al_6076534a,al_a5f7e6c[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7e31f5b3 (
    .a(al_7b59c46e[31]),
    .b(1'b0),
    .c(al_6076534a),
    .o({open_n109,al_a5f7e6c[32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a7b3404 (
    .a(al_7b59c46e[1]),
    .b(al_f12834e3[2]),
    .c(al_dfe2f2a3),
    .o({al_dbe911b7,al_a5f7e6c[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e8fd128 (
    .a(al_7b59c46e[2]),
    .b(al_f12834e3[3]),
    .c(al_dbe911b7),
    .o({al_a7fbaeb,al_a5f7e6c[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b35a80f6 (
    .a(al_7b59c46e[3]),
    .b(al_f12834e3[4]),
    .c(al_a7fbaeb),
    .o({al_59bca917,al_a5f7e6c[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3af992e9 (
    .a(al_7b59c46e[4]),
    .b(al_f12834e3[5]),
    .c(al_59bca917),
    .o({al_c92e4639,al_a5f7e6c[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9744ace0 (
    .a(al_7b59c46e[5]),
    .b(al_f12834e3[6]),
    .c(al_c92e4639),
    .o({al_a5d442e7,al_a5f7e6c[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4f418d2d (
    .a(al_7b59c46e[6]),
    .b(al_f12834e3[7]),
    .c(al_a5d442e7),
    .o({al_91974942,al_a5f7e6c[7]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*~C*~B*~A)"),
    .INIT(64'h0000000000000100))
    al_78d54170 (
    .a(al_25fbce42[5]),
    .b(al_25fbce42[6]),
    .c(al_25fbce42[7]),
    .d(al_25fbce42[64]),
    .e(al_8a4a038[5]),
    .f(al_8a4a038[6]),
    .o(al_f036124a));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_3d2fbb21 (
    .a(al_25fbce42[4]),
    .b(al_8a4a038[0]),
    .c(al_8a4a038[1]),
    .d(al_8a4a038[2]),
    .e(al_8a4a038[3]),
    .f(al_8a4a038[4]),
    .o(al_6291136b));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_5ce08aa1 (
    .a(al_f036124a),
    .b(al_6291136b),
    .c(al_a7af1013),
    .d(al_25fbce42[3]),
    .e(al_8a4a038[7]),
    .o(al_a27f756f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(C)*D*~(E)*~((F*B))+A*~(C)*D*~(E)*~((F*B))+~(A)*C*D*~(E)*~((F*B))+~(A)*C*~(D)*E*~((F*B))+A*C*~(D)*E*~((F*B))+~(A)*C*D*E*~((F*B))+A*C*D*E*~((F*B))+~(A)*~(C)*~(D)*~(E)*(F*B)+A*~(C)*~(D)*~(E)*(F*B)+~(A)*~(C)*D*~(E)*(F*B)+A*~(C)*D*~(E)*(F*B)+~(A)*C*D*~(E)*(F*B)+~(A)*C*~(D)*E*(F*B)+A*C*~(D)*E*(F*B)+~(A)*C*D*E*(F*B)+A*C*D*E*(F*B))"),
    .INIT(64'hf0f05f0cf0f05f00))
    al_9ba132d7 (
    .a(al_a7b01c14[2]),
    .b(al_a27f756f),
    .c(al_5c72a609[0]),
    .d(al_5c72a609[1]),
    .e(al_5c72a609[2]),
    .f(al_25fbce42[2]),
    .o(al_74dc1091[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*C*~((~D*B))+A*C*~((~D*B))+~(A)*~(C)*(~D*B)+A*~(C)*(~D*B)+~(A)*C*(~D*B))"),
    .INIT(16'hf07c))
    al_76443ad (
    .a(al_a7b01c14[2]),
    .b(al_5c72a609[0]),
    .c(al_5c72a609[1]),
    .d(al_5c72a609[2]),
    .o(al_74dc1091[1]));
  AL_MAP_LUT4 #(
    .EQN("(A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfc80))
    al_e7514b14 (
    .a(al_a7b01c14[2]),
    .b(al_5c72a609[0]),
    .c(al_5c72a609[1]),
    .d(al_5c72a609[2]),
    .o(al_74dc1091[2]));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*B)*~((E*~A))*~(D)+~(C*B)*(E*~A)*~(D)+~(~(C*B))*(E*~A)*D+~(C*B)*(E*~A)*D)"),
    .INIT(32'haac0ffc0))
    al_a1af4d2c (
    .a(al_cb807890),
    .b(al_6380dbe7),
    .c(al_e7b5abb5),
    .d(al_a7af1013),
    .e(al_4fc7a4fd),
    .o(al_8d6e0488));
  AL_DFF_X al_29fafda3 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8d6e0488),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a7af1013));
  AL_MAP_LUT5 #(
    .EQN("(E*A*~(D*~C*~B))"),
    .INIT(32'ha8aa0000))
    al_8e2c06ab (
    .a(al_a27f756f),
    .b(al_5c72a609[0]),
    .c(al_5c72a609[1]),
    .d(al_5c72a609[2]),
    .e(al_25fbce42[2]),
    .o(al_cb807890));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~A*~(E*D*C)))"),
    .INIT(32'hc8888888))
    al_40419603 (
    .a(al_6380dbe7),
    .b(al_e7b5abb5),
    .c(al_fe97bdd9[0]),
    .d(al_fe97bdd9[1]),
    .e(al_fe97bdd9[2]),
    .o(al_6d2e3f3));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~((C*~A))*~(D)+~B*(C*~A)*~(D)+~(~B)*(C*~A)*D+~B*(C*~A)*D)"),
    .INIT(16'hafcc))
    al_c3f2981f (
    .a(al_cb807890),
    .b(al_6d2e3f3),
    .c(al_a7af1013),
    .d(al_4fc7a4fd),
    .o(al_3660546c));
  AL_DFF_X al_2adbd347 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_3660546c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fc7a4fd));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_d7c13a9b (
    .a(al_b799bc04),
    .b(al_d4a46bf1),
    .c(al_43722bf9[0]),
    .o(al_daece8d7[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_570e7e82 (
    .a(al_6893b11d),
    .b(al_d4a46bf1),
    .c(al_43722bf9[1]),
    .o(al_daece8d7[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_825693d8 (
    .a(al_52c6af0a),
    .b(al_d4a46bf1),
    .c(al_43722bf9[2]),
    .o(al_daece8d7[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_3ce67d3f (
    .a(al_6f63d541),
    .b(al_d4a46bf1),
    .c(al_43722bf9[3]),
    .o(al_daece8d7[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_217c2cce (
    .a(al_69807e37),
    .b(al_d4a46bf1),
    .c(al_43722bf9[4]),
    .o(al_daece8d7[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_eacdcf8 (
    .a(al_e7b5abb5),
    .b(al_4fc7a4fd),
    .o(al_38acf7c0));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_8891b6f7 (
    .a(al_e7b5abb5),
    .b(al_4fc7a4fd),
    .o(al_8143d2fb));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h7304))
    al_a616175c (
    .a(al_6380dbe7),
    .b(al_e7b5abb5),
    .c(al_4fc7a4fd),
    .d(al_fe97bdd9[0]),
    .o(al_6f31a76));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*(D*~C)*~(E)+~(A)*~(B)*~((D*~C))*E+A*~(B)*~((D*~C))*E+~(A)*B*~((D*~C))*E+~(A)*~(B)*(D*~C)*E+A*~(B)*(D*~C)*E)"),
    .INIT(32'h73770400))
    al_3742b29b (
    .a(al_6380dbe7),
    .b(al_e7b5abb5),
    .c(al_4fc7a4fd),
    .d(al_fe97bdd9[0]),
    .e(al_fe97bdd9[1]),
    .o(al_c5966d4f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*(E*D*~C)*~(F)+~(A)*~(B)*~((E*D*~C))*F+A*~(B)*~((E*D*~C))*F+~(A)*B*~((E*D*~C))*F+~(A)*~(B)*(E*D*~C)*F+A*~(B)*(E*D*~C)*F)"),
    .INIT(64'h7377777704000000))
    al_9d303a8c (
    .a(al_6380dbe7),
    .b(al_e7b5abb5),
    .c(al_4fc7a4fd),
    .d(al_fe97bdd9[0]),
    .e(al_fe97bdd9[1]),
    .f(al_fe97bdd9[2]),
    .o(al_e9ef2594));
  AL_DFF_X al_26b40ed8 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_6f31a76),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe97bdd9[0]));
  AL_DFF_X al_4ae1a92a (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c5966d4f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe97bdd9[1]));
  AL_DFF_X al_65e9dd52 (
    .ar(POR_RST_i),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_e9ef2594),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe97bdd9[2]));
  AL_DFF_X al_933064d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[9]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[8]));
  AL_DFF_X al_6e5ee8d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[10]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[9]));
  AL_DFF_X al_558913 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[11]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[10]));
  AL_DFF_X al_766d3233 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[12]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[11]));
  AL_DFF_X al_caed43b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[13]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[12]));
  AL_DFF_X al_cf1a7ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[14]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[13]));
  AL_DFF_X al_abdd07b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[15]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[14]));
  AL_DFF_X al_bb51d58b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[16]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[15]));
  AL_DFF_X al_a5556141 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[17]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[16]));
  AL_DFF_X al_43d89ec2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[18]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[17]));
  AL_DFF_X al_df53abb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[19]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[18]));
  AL_DFF_X al_ac43ca30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[20]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[19]));
  AL_DFF_X al_1f8bc185 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[21]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[20]));
  AL_DFF_X al_3efe9cac (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[22]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[21]));
  AL_DFF_X al_3998118a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[23]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[22]));
  AL_DFF_X al_d838c1cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[24]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[23]));
  AL_DFF_X al_6bbaeae (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[25]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[24]));
  AL_DFF_X al_1d36ff2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[26]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[25]));
  AL_DFF_X al_cdf220c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[27]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[26]));
  AL_DFF_X al_c8491c4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[28]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[27]));
  AL_DFF_X al_b5f73a84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[29]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[28]));
  AL_DFF_X al_c7e082af (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[30]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[29]));
  AL_DFF_X al_dfc6f8c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[31]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[30]));
  AL_DFF_X al_27c4c541 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[32]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[31]));
  AL_DFF_X al_1f4378e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[33]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[32]));
  AL_DFF_X al_651fd12f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[34]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[33]));
  AL_DFF_X al_4a97865c (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[35]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[34]));
  AL_DFF_X al_9dc7004a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[36]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[35]));
  AL_DFF_X al_94b0cfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[37]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[36]));
  AL_DFF_X al_78859365 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[38]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[37]));
  AL_DFF_X al_e8c96814 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[3]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[2]));
  AL_DFF_X al_2449f65b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[39]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[38]));
  AL_DFF_X al_8f42f62b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[40]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[39]));
  AL_DFF_X al_219141d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[41]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[40]));
  AL_DFF_X al_39b85e30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[42]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[41]));
  AL_DFF_X al_99c7484f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[43]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[42]));
  AL_DFF_X al_a388632b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[44]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[43]));
  AL_DFF_X al_852b84f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[45]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[44]));
  AL_DFF_X al_d4be563a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[46]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[45]));
  AL_DFF_X al_6db10125 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[47]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[46]));
  AL_DFF_X al_52ba6f40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[48]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[47]));
  AL_DFF_X al_93cf1c51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[4]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[3]));
  AL_DFF_X al_30f761df (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[49]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[48]));
  AL_DFF_X al_2d9d65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[50]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[49]));
  AL_DFF_X al_727d1106 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[51]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[50]));
  AL_DFF_X al_6448bd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[52]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[51]));
  AL_DFF_X al_7f673942 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[53]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[52]));
  AL_DFF_X al_56756846 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[54]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[53]));
  AL_DFF_X al_2b9be308 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[55]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[54]));
  AL_DFF_X al_b2f8d39e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[56]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[55]));
  AL_DFF_X al_8dd20261 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[57]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[56]));
  AL_DFF_X al_53cde693 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[58]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[57]));
  AL_DFF_X al_f1d6355a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[5]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[4]));
  AL_DFF_X al_a8a8934a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[59]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[58]));
  AL_DFF_X al_ac039c82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[60]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[59]));
  AL_DFF_X al_d878c66e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[61]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[60]));
  AL_DFF_X al_c6fb719f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[62]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[61]));
  AL_DFF_X al_4ecd660e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[63]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[62]));
  AL_DFF_X al_5a4e5f73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[64]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[63]));
  AL_DFF_X al_85941634 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[65]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[64]));
  AL_DFF_X al_caf01a55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[66]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[65]));
  AL_DFF_X al_a5759452 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c2ae0151),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[66]));
  AL_DFF_X al_29a1237f (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[6]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[5]));
  AL_DFF_X al_c3f655b (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[7]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[6]));
  AL_DFF_X al_c4b5c385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_25fbce42[8]),
    .en(al_8143d2fb),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbce42[7]));
  AL_DFF_X al_5f109b35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8a4a038[1]),
    .en(al_38acf7c0),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a4a038[0]));
  AL_DFF_X al_b9acb776 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8a4a038[2]),
    .en(al_38acf7c0),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a4a038[1]));
  AL_DFF_X al_a7abe470 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8a4a038[3]),
    .en(al_38acf7c0),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a4a038[2]));
  AL_DFF_X al_52469b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8a4a038[4]),
    .en(al_38acf7c0),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a4a038[3]));
  AL_DFF_X al_a2bce94e (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8a4a038[5]),
    .en(al_38acf7c0),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a4a038[4]));
  AL_DFF_X al_a0ee6413 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8a4a038[6]),
    .en(al_38acf7c0),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a4a038[5]));
  AL_DFF_X al_7ce74c0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_8a4a038[7]),
    .en(al_38acf7c0),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a4a038[6]));
  AL_DFF_X al_75126078 (
    .ar(1'b0),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_c2ae0151),
    .en(al_38acf7c0),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8a4a038[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    al_3fdd5e3d (
    .a(al_a25a6119),
    .b(al_fa66b6a3),
    .c(al_f0ecd262),
    .o(al_3f2c3141));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_8b87d4c5 (
    .a(al_6499e5fd),
    .o(al_99763382));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_721b885 (
    .a(al_1a1af7e4),
    .b(al_bb0cd305),
    .c(al_501dbbdf),
    .o(al_a96ccffb));
  AL_DFF_X al_731d1aca (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_a96ccffb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0a7a5f));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_a96a1821 (
    .a(POR_RST_i),
    .b(al_50debbc6),
    .o(SYS_RST_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    al_11e57a7b (
    .a(al_1a09507b),
    .b(al_b8fe1a1f),
    .c(dBusAhb_HWRITE),
    .o(dBusAhb_HTRANS[1]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_5166f2a4 (
    .a(al_ece70a8c),
    .o(dBusAhb_SEL));
  AL_DFF_X al_8eafbaa3 (
    .ar(SYS_RST_o),
    .as(1'b0),
    .clk(SYS_CLK),
    .d(al_afa99249),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aabf3e05));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_fd73cad4 (
    .a(al_ece70a8c),
    .b(dBusAhb_HREADY_IN),
    .o(al_afa99249));

endmodule 

module AL_BUFKEEP
  (
  i,
  o
  );

  input i;
  output o;

  parameter KEEP = "OUT";

  buf al_650f98eb (o, i);

endmodule 

