



module mipi_dphy_rx_ph1a_mipiio_wrapper #(
    parameter LANE_NUM = 4,
    parameter BYTE_NUM = 1
    )(
    input wire                             I_lp_clk,
    input wire                             I_rst,

    input wire[8:0]                        I_clk_lane_in_delay,
    input wire[8:0]                        I_data_lane0_in_delay,
    input wire[8:0]                        I_data_lane1_in_delay,
    input wire[8:0]                        I_data_lane2_in_delay,
    input wire[8:0]                        I_data_lane3_in_delay,

    input wire[LANE_NUM-1 : 0]             I_lane_invert,

    output wire                            O_hs_rx_clk,
    output wire                            O_hs_rx_valid,
    output wire[LANE_NUM*BYTE_NUM*8-1 : 0] O_hs_rx_data,

    output wire                            O_lp_rx_lane0_p,
    output wire                            O_lp_rx_lane0_n,

    input wire                             I_lp_tx_en,
    input wire                             I_lp_tx_lane0_p,
    input wire                             I_lp_tx_lane0_n,

    output wire[LANE_NUM-1 : 0]            O_lane_error
);


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-009"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
atMwpWETLBZaKKSJbBuPvE9O7jvKhFlg5XqFNyixWGX7oYFwZoa3Zte+hA3PS66Q
J+KkcohxjO0GrmvPyKMf5ptPeBvNfZVxJF21lKVQKi9mqCg9D47akqGKMMsDCzk/
GtAjoIN8zx8qJhtFVMgewepFmV8TptbaSUSoabhPDfU=
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
A1SuazA57hiGZQdublEZ9ni2nv3q6F5V0OBO1WSKt8ddUX/Rd9TkBtO4vt4w04Dk
HQNw6sC5RBmLL44eGBVQT1XtoFEuIWpA+VBQMgoQ8ie98WhMtos06rpZKR0GXJoI
gcLZyXqazaE8krOExQSA06tJiKZlZehBXxYuffHxPc9h1IMsUwBy3ewcP6ptyxzc
zdrkN9Kx1vLtCysy6hHHMq/rVYKjh7OHGGSVcN1QVKgO8nYHjbhBVbFTUAYb2MAJ
Zr9lUGame3hTSIh/P5aeCfmqQuHqOuzkQ9TL0YEyzHgtXc2H4V18fhHEXx3b+R/H
L65MJjUTGu2rrFz1a18L0w==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
QMJ3NMcGYDJOL91K3oGsdYfTOM2W6I9ww3MR+E0P8VCgsXKrJFM4HdBgtPKbKATX
yy6fMhmL1reUkbGSemydIsUnMXWJB6/OhH48HpYFuGBkBSVauGoMcqC3iUyi9W2m
kswt3rAATv4dSRQAjlzFpyU2195dOlrtRWSEO4k8ZoM=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
YJep2igG3zJ0f23RIbPlsDz5Ih+pQOWfnyVvRkHkcisBgQS04+IqUkt9i+/WLwTZ
E/2ZKNAqxgGydy85o837HS7LW0pcYe9nTWnx+OL2hbpLwBgfsYZNxpL/1xxPq7lU
QEqi9OeO6CfMsrx/xi2XGvhfIUF6Pq1XDkJ22UhcnjbzbiZn8CUUndkk1FKpM0ve
LXWP9NJ1dlFUkr1qyWzqVT1bD1TqgpVhGW6KrqZrLaM0kY1fMSQhF5C+IUAMuQep
Y50WWB/Ps7iG1kCagW64/p0xbzvDte8eYSuvyb3Y0o7n+FeADt7P+YpvgS8weCSS
O3dqotTIKm0Nl01vnF5gfw==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
PmDVEH6sHG7goSIzj1eaEUuLJ6ymaK2Mw0tAswUAJXv/u7raxblM4YApsIgkA6qy
a3MlrFy4SJsBiHrEVJ4Sgj3d4lkj8a1VpZ97A54SB4tD/LRtUCWcvjN56i0y/Xzg
FamCyJEOLJJX9x90tpFVw8S6VWyEUCasLmDpHTK1MGg=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 40672)
`pragma protect data_block
5lXjm33GM8xpKhLBd7Fx1RY8jvTIRs60OofZqyiZZuEQg8c+dt62u0ResKXoenZW
3hFvPuKngMoZRgwrN+gam/QWRD9wMwvkXFuQuemKHtmOpx3zim8pyp+v5jJynNkB
lus+AfdBv8QD+E7wWhz7ZzGXdEzHkyErOj7qHa/bD+Y9SAWftaOMuPKUCeBMeAxE
yzfT2cQpjDNcckDxDYunymBaVA4T7iqOmoRME/0Nyas9q275LTXxrQNvXZmaGMT0
285On1rMGWrtARutBxmtZuvuI+SnGjdZJCaQKl30Rkly1Jztwlwbo+uPyIpQwV1z
qnD0bfKtkg5/sFPmizSArqOyHBGjk6BcBbi09idMh2b7y3tJiOzZlyckXS5XYEad
IWedwdScKU3q8t3pYIGFTTQr8qrQRYd7Xq0elQWfaUAjv6X7YZpx/duNDtnmORR+
0IItlHOe4b4L1Mwvl0mynGz7v2Zxxsodw8FhxARPca9Efp8jz89VY8SgJ1Jim1py
8bgqVPQQA+Swwiu81kW0vuRr4QwOxME2tLMyMPb7hzq1SN+cpY4V06zc7aQvImDM
nGcW4kcyK5ZfWaaPE6Q1v4i+PyEah4X9W5W52xdb3UZdBTMIDPRUubYhv16XHz/4
esbIh9ihFjAph2q5VrwhpHZ3e11ekmvadFLAwDmvMaD6isbnjcD6p8ZWuftq9GJk
CumFbCCcWB0XjKi3tXN0z0ueJD9Vqztrqbqbs+MOvv99LMgwxtyCi8QWd8W58C8D
9TFHITQT8WcSjwXbrotBQDK6qkCEUWd5nbx9wO5r1TTPnsTukPvbWmAmjDVX1xUU
bhCtzn8WNMWbUJDOR+4mH0iThxr0YDTn8rmd/SiNzJH7ZyVvSnTUbU4adQ++sDiQ
Mhv+bOz9OuK7A4Z5YYBnCFkhQizJm/2OVHWzJvIFQAbnhEUiZCqT7ghYDvc+E+Cg
iAXFP3IG5EKyIaKc2EEwjR46s+AnDR+BgRYkeMIAhJuEH+IDxNgeimZhx7hCfuCE
ZBbJZlfGKm8DKRs95emRqPBxCpLScyfN9YdWtYcN6faOJsqyp6LYG3XZpX66Zdvz
xMl1XLyXL0I7DAWGOzQHynTgAi8orxCAgdu54jOWj4ytKiwLzEFA7r5CAHXI5WkC
C6dGSYgufhS45/JMCok5gSObWbEUcosn77FA2bbPv8G9Khb1MPuNU+1rpdo4pbXM
U4udi1LpgsQA3qeGB2NvbHbD6jHAo4GdOfY8jRO1fgwWUlZSW4ZtBqrfKJiRB+rK
KTDM2wSSL2AZ2x28oaMUSn5sVbLbMAPpZSkYGjdJZkxZ8Bs1AMU1DLiZ6XWEwYSb
PEyaUk442zcWE4aEMj7zu8F2nTs29DDeaTozakf/ku0VeVFdCGA8oFa10QcIUyuX
kCxxO2jWSqDurN2gGfreRbP3ygrwP7VP4Zr6vNBtAtvFJ93cy2bvym5up2Dn0+f9
yDXqzi+L9U8tbXKC1o+inD6x6vY7j8j1mP4W5Bti89zKGgRXoQ120PMGM6UpM9e0
Rn6wnUrIyUwbEKe2hekv8p6f0n2bt42258ZfBHQqizZvGd/0ygD4C+TZz9w5S0b6
ln/d8943zD+7qKFxDghOa6Xq+pFChiSVb171LAWixiJEiNYoO9nV6OA0Rd1Q/iKW
NKc5w1NIv6mdxMQ0IKgLyUcXnFGSdxXB2XSaPEG8kUkmG9JX9b4Fj29zPiCQ31XG
DN4oWTDS/mJJYjSAgHy5OmuBtQ1iyoM6dy0jjYePTzrEIRsM3s8Lyx5ZP/KwecKs
nated8HtGyodCEHy6jsrfOIWXL4CrbVGrk+71xqbYlsO1QulKlFlfdHdKzY60cDn
4mgY1Cq8d2rBWD2z+Q17nLC627i7XggtrvjnnavhB1OZRWkGDb6pOaEJ8Xdtntct
VI1FSKIJZqxwFNHT1UWsUUIWyW9JHaY/T3oeAWBtbxgoE3yLA9djOjo1r5hZ0TL9
eHqk+V8O771V/YTNqcwfWs7fKDOdj2vTGfDyUb5T6vCFaAVF6lTnsHr3IbR2RKmJ
woLR0T269cv8VzpJxEugFTqMQ6SRo1cfKkmiSlNyw+aURP29jvFCJD3cbQ/3dgLZ
rNO8Gp69GJG7jVeD65TlIljfBpt58PFI5so1y7P31VEfCGwa/c9jLqd2jBFRwm88
rkra94tKvVHYxVgoqzfd9SnLjX8PNaqcAwTR9Cd/Ai0UfeWvvlyBRFKX+p/aGdaX
xRGjFcbVLfpPwQGJ/CVvdikBuJ7jmggWW0cdcZ3kTjhP1QluNOfjMmOiO+HDwbx6
oBihSGfWGcDL/WdDN88sBpkS1NhVwWxuAkDXXXKy0UuJ+0Akd8iN6Nrd5ifBVXU5
OzATmoqScZRNXZ39+q8StPp8rY1N1vuQAyNoWRHujWKcG3Uu0hDxJg4Mn+delGtj
ADWAT+MxBw67oXBEG1e/r9b9xvH5yvCTGIyAp3+L0fnL+eLfcc+7AOqf+dc3Y5/j
HQI/W0oTBTJd+cSD3Od61jG044FAsWg1xAQXRpjsx2ffSfO5qeOqsjpQctdBH3up
vJEuIPrp5+jqlkPmuLcNC17P6LS3SS7PuSqFHRcdJs/ZT76x4FVk2vRIRfAbLzWn
gnDITK1cuyL6EP68OnSWQsTcj0SDtYrb2mALV8pYVlyhrlgajnoQOhQMjwo7/w06
ubRu1HjFb8t9OeNsuqdRUrFM25aRE2GR1Ix3vz4Iy7ySeCmaEVMayFxNVsQcwiOm
cHMGqmi7zO3Sho6a2go+PunjEyffZAxeqGq9CUR6GY7X7kW0p4mUrDYONOd3P75R
dEOe6jDFcoeZDzKzUK9fqq4VCcf0HbeqV8F8ONFfYWKZZoby3GqzNRMP4CXo75JH
7pG/I7Nzr9neNmf38T35MxYFJtfugOvjxYRqox1nsjBsKT9issgNzYDHJv3Bhka5
zdJ0juT7IuyThKGK0yUJI5u5pNt8wLbIbujBAbfbJVo2eZR6ixFGNs/Vp5UPHOJZ
JUc7fbUjJtq+r2NL5HxXbNi/6HEndpz3xLL/AdoVmWW4d9MIugqxyIzVB1PCcaeh
qO+2PKLM585j6b0vvASrQCtcny2PDawMGR40j0OBBuIWQ9Ep+lP5ochE57U8MsjE
G6JchMKxa8jV2YSftyy8Di1g3kygR41mngtL9nzwPv5k3RD2IENhLZE85j9XF+RB
D7lEeJCxyHW4b5vYTyhIMhjdFXVNiADHF8EAVZ/A5hPqVEMVIFRCVpdpSuc7b44K
HMlQOB8aBj/ahYw6P0s5p1w4M/xPJuFfomO8+jLKOc7jPFGJcvfbLxNZq2LJWyMf
L7Cca3MzRNUPK5sK75ciLH7Tv0Bi6yOAsTzFg7UnPmSrhP8TRE9CU/JrHAPfsvzt
e194gOpawSuEk9xO3UHE7OfCYjUcR1g0vEVMzKnotjFL+Ifldvk5wZBX7aR1Au6F
IY9BxGL2deWiTjbXWH9GfhNik87ymnV65OLXjK13AKtjwWAZ70RLak43xe2dUNN6
nfqupo6lwq4ji+SmxLJnR20gX8apkVG8UzRAwQJBeFeaBRdRV4a0mVMsaQAmx5K+
Zhz6OX+bZuD0M7cnR5UpCcgbMRe2UOctiCS4/4HWiSR460Nh35P6Gra+8Bmb77Sq
xHtOhA3eEkholcuwyGEhJpNViT+HCOtibDJoM7vHB9ETHq4nY7u3Bfdcs4r9bJb9
wkxNLQKuWGbRJnhiIVODivyhC/fG9Lq6/DSIeERgAgEac9xpzJU1JdAsqNR6OQv5
jAcm7LpfcV7o7Ha8R58EIUZLH6Wmy29CZAejIBhQe9Hc0RYJm/pYD8mjh9LMg+Dz
IxpE0J3gPpT+A/ptKnxdNf1m83lFAhXgF1cXs21wPP2cHSq1UCorILsKizaJ5M+A
/cD74L+LvIgNczbSNPK3wmdLMoI1WC1GNZjyXkPRJLpU88wFDVZdvhj65pyx37Ln
teUjWewyvMPP0IHjELLQehjPkNdNy1tQHoygA0/5oTJel1B3wjXJlmm6pu940tzm
5IRgLAmdERxgFAXFTbROE+hjewKkq8pNnY0wBTPdtaQKyaPi5QD9zoeeMzE+xCD3
O30gIOJIfrs04sEBBuunUd5qpqd2Fr/DQtXqRcPQHxwoPZOP0T1E116/f1g0Ld2p
g0lW9OitnShl/c9PteKSivbmIIOTlr+LaTj5twj2jrM+z7Wb/isT3zKRqvGpUGTC
PJiBtebvi00DA7+3VAKZqYDOjsAJnXb+5H2L9h1Who2PgzE2y07uOkPZymx5U8/I
FLP+Da9X8uXHazm7Ma5xWl0U5TD0IJ1N3fryqUA83NdcuF5pooeF6+IKtfbPCsLh
sO6uA6sFgRml+X1FnJLJowmYG5hLL73p2Xm5HuQFeCsDk1u6wtlWI9HrRpYf6N4C
LHjkot0ngh1b1QPRnsOPO6pu8+bCn63m/RXk+Fk/acULTjusPlGVjUOa4T4xzIMo
5c4HJU0n6BvGF/dk20b+mtiGL42uB42OuS/V5XgNtzi3rwMFoQC9mXT1KQSAmogG
zq8ODUwrdcacSwO8y8ozrGNE3UwCMJHQ8UqYz3dczc2g0pE5QWLK4RT3L8uwZAgq
Fxi8aMkQSF7+n2PjxjmNF41jAHMnIJLMeRGt8ZXtHJvMTbuO3GqV2abc5BTHc2fu
OOTH57Y6UpU39p92sbXc2pGjiwoqhTTz6oRTgOXMYsG08hKf/CfW4geg0QyVBZPV
EXFqnEBPA2aeCvNPhY/98kJK8CzkK3trbjfjIHlwRwhKoG17z5nZgNBzredwfJze
7pMJZWCQBrhx+o6ZOv8b+pstIcIhUqRib6wF/pKtBSdkGiYL5pyN5EnOJw/AgkU1
qnS4tp0ZXZdvyAoekQc/SEmdLa2f1ey6UQOM01ig2EnYd0lxuBASXF/y4wK62FEZ
IdUWjc0O3Z+MqzJiN4Pb2jPHokNtjxM2jPQ55ERw21u8BUhUplSWnuEzPFozv+7/
auNHCYXAIY7Il+QM9tJotXu7te0xHsKwKVb8sN/+jF6tjlIXcoKt6NC/brWUV8S5
yP2r/GZ+zF5pwgHlmXGKiJCYV5PnIiuxT91Mzlk+nSEsyORnB+tbOLleqZoocjdN
7UQmY5F0hf5UjseyZ5Gn3gLB2GREWqlTHnaMg1QjOJQlPNb3dTNwGdGRxS3WIoAX
XQ5IqP3C/kbXWZGOCkQq5KtFdZuzzoz0nlPbNelkrJuvYb6zHAdRaPEE1ao/irwD
M6xsfrtkOhmeWo78RZB/eF21+hKbtjWdL1D1wv26kvpvAVQJdaRa0t4V39zfiGq1
Q8cbBuBGQI3GnhbX2IL8h6eUg3qy9sCNHgKYwwugkUj2vwInHOJMiNbgH2okwLGs
MN2X0aO96htAwef8Lu31BVPXM90wAFt9yGme6adtT4a3bFjMSvKgHyX4H4T7BfMx
ySnC1YxKNZAICvdh/SysOwdSWiIRdV0yZ239U6dU1rAsO8URzOvWSKCYFfbCnny3
a7600X2lXRAT3IRUtMlJF071Fp3Sbav+/eqTn6/UcjkaLBIZDVBt5qKEWeYrYBz3
++3rymwC8TXZMeIX59oxPKjK6XGCWJKcOYXjxImAWkcuLpqQCIq3Uxr+bbLi0u4w
TRIU4ok4KB04YHT9eduDZP6q1foh1BxJ3yeAjfB0XpEOznCdaBX4/exuAPCoaY0u
/HBMw1qsVfXCFkBBjLVW33Zbq6Qzs1ziJAMzhesZvH/sF/x36nfI7bclEzxHjlQi
/4spzjk/0n7l6lNmAq9j8+kWMGK8mXgVrWwHvyvGxV+X9tNTdQrornp0470yzahi
rjcYO+y3GZ4z1LHY663qf3HrszUeEfeBZGpHYA0p4zISRmseeqnTh7F+2ID4/DSR
QdmVIjRtXE5Ce3Ot56+cwdFx6Png6W4GSSrm3bro/Z5hWZO8o/qiIfvXy6HSNi+M
UZ/j1XqGxMhXcdz1h6/r0ZSIMFFEHWk3liF4LiE+BU5Pb+tHTnWpTjElIFEYY9V3
4V03nKXCebevni398tX8zvZNLNNU7CNq7+mU7DDgipoaoWeee/iHeRf8HcImKHGm
s26pWNI3IFV6MV/VHSsK08LPYwFgkoaWCQbEdGKV4gfbVEOgMur43nmf/AjFv6fy
OQWOYT6DrFNOSKNE33zsEEuIm87nUjf9kuTr7Xtqo0sF4XglmBt4l+dyF1FExPEP
UiNAVMb3tf+96964+suq0SvBEWC79+N99rxZVLDGoq69/prHsnQZh24eLBKHGB1E
UROXFnezBLdM05+tfny9zewAiJmoTooNsmFJhgaPohHJ0B8FQOzwz40/VkqjV767
Fo1RHIBzoZdVbAonkMBHf5oqqDqZ15ejsfIWCfgliBbW0qR41ENqwSgDZWbo5Ccc
hpfZO5yTo+2v3xU/tBGMt3SqZVXChFlYeP4f0quUGMo/qBLWwUtyEmADxsD9bPE8
2y0PAFEs6kVaz8wJamx5KMkxRNsjVX5sNq8UdBaTSBqVeEGMXNoyR3OkA6GnJ89d
wGP/Et5ue0rYktPLyeZIMRQEHgQwbTl8SPM9osbjMe/a3W9y5UwsiTOWjthhol+k
7bY0osv5hp0SdsZOva7rhx9eRpPmKP+bPH5imhhYz38qEr5uywjJlxm/LvuwtHKg
EaFDp0N5Jk2gmcOqJmosmfoWz+tVySEbm6phn24/D5/vpObNlrypzQOf4cEGxmKB
6xAO0niYBYxBPJdx66cHGffCkewRNOE+2l9lho7yI/x8nK06xXocUIfJOWuBcZVf
s0LchHIokIUCT+aM2lbBkQlYaTU8pPxYvNw8EBTJXpHxDcP27JVEsoVJ7baRvvE3
/bQGV+VMUxmBI7meaY8Sw3I/iJsoslxWvHHD69rk5ZmVWLaF5efp5ZWy8b+7kf3F
Ova0kDIkC8T9ukwF1YeYMYtjG+JXQZoy1OV8bFxGjuarC+CsJUYVH5pIFglYzT6b
2M6RUpf3Z3Ityd3oqGHuah5LRmVVRHUNdLT9A41EhsY0gECDTUC88gclEBPDnE3O
ua0lEdxvutO8Qa7Ap4xv2nVaOZUi9Btz+Wr9iyIdCAHi+oC4puAdqCEkEbmHbZWi
TOWaEKxL7eIRY35g7owm4BBjmH31klcmTvCb8b1At3cI9bg1Aw8fO2Lm/00s/en6
r/ahJ34zX6+JAZz8rrAL8MFc0c8M+helPQL5pSQzp5iKHiZ+ubiV7CnwwwNChGlY
Arle6Sl6f2+JookgksgfvWEKC2Nwf2zzYIydhrC9GfV2SZ6ASTmJMvyqgygAXvTB
hHnCFI2G4XWvcauAZvqAiulflHGy1Qw2ALvp/7CZJYOSHsqSrr7nDGj99jgS/IHM
PFqmPFfUjv49E2Ht9qgw9Q1LdayjzMeaGBYbBzMLrNW16IdOtBTt3k+0SEqCKEaW
Hx8fPMFUKugmX49D6mBKwJti4LCjq4K+mgHpat9HvMv2qrs43UV+hzsa7oLeTo38
XncplG6YdhFRu2Z/zrWAc00HRKJwF/BUQAJjaVsKE92fy3DP5LUGwUaSaji/T1Ez
RRGGIHLP+erOfEyPNgR57fAtubIKoT6t6nNm0DTVouaCAjf+jl3TCdS69WDSL+D/
UfEt/IyPyc0Q1tniCzH2IBXuRU2wtvMcrVgsFCeeYDHRJL1jM413ankZtE8635PF
1kRfbtFm/s6SJ9NtM73ggMik+68IfEEaNBIrD8PALAj2Be9PGqFC3mX6nFz1V/9c
lqurPQ4qV6I7ddKT21qb1d66eNlAfBe9uUN3/HvHN/9H860qNoLtLi20nMjzZtvp
J3dqDaUpAJ6LVJr2mz+nCo9S/4dODmM0idntkCdEM81Y/5OnvnkurvVMRHo3ySrs
QQR/QdCnKFGjpGa55uJI+fM6qV6r9hFmfM1d5uhlKvMY8tpH0kBfNdgNLAa11QrV
QjejQN8/1YbXSG5zOh114rJcw601e/PG1FuE3vNg5ayS1d5v3elpeTH5XVfLgcnJ
bbBBwpWJkl8bKHPXSKK7N9hDup8e6J1cr/IPP+Li7ecYki1hXfpw0lj5hctH48Vx
Ld0HZH+/UnnIwI+I84uU6jGZoHnJRGNzsiHMI2t6KwyuGjFovQgo7MCQqo3bYGUD
vvjI7DBUnEhnH5WJxkdzvm7msmX5M+Gebl4JqpnrKsS/5MAerp0N+lZKEwjxe5ZV
tMceAUCyxgdg+m5zVqka+m83DbDKMIo3iZ5tC/GhpWQntIAJdHtE8OeX4v3JtAdK
obxHudZ4Mh8FqPIG1rnQgPG1svI+it0ANTN74lMZc8cYqavxv51XgSAHB7BD8Ug8
CNtnb6JxN77ZSviHmvVS62Acw/ypU56lxb+EmPUUozdRozXVKGHZ5c9XAb09tpBC
bZC1Aj485iVbVWlQGHZbFTIZHRUOZj7RfjxCmQPIDXVy9n3Jdb5OuBeQpSL0yx4C
aiwNOo3X118aX3dvgCWYTzxlZUU1mjZTnAD0zfgymAippagXeetItZa2q/ddhUf2
N4OHtQg905Y7i7yC5KNKe3lyAoDmBQB/rP+bydgIIiOj9YPOGugWW8O9vK6wKYJK
W40hA84wd/nDMYuKzRKoYWsAYCvJXO2UPFQyYUqqsDvbGApY3Kxlz4o4BeH3dBXi
3gOCekUNN20R2pkPYEZY5YuTrucUveL/EugX43YJM3Ltop16S39KBrU3Uwgf8DcN
qlw1jcdxcSQ+kTw3fGh4tAv23kBtbVOi4NTCqVZv5VK7ZLqDP+YyOvnj9TPdizUN
VeegqGt3yMDdD5VmgGRtkDgLQTg/XvSm6yqABmDeTv5mbFjt3V6kINwc13eHAqOr
2BuqTZEXNrkyweJzlzvdhVBR5XhH8pPhBcyw/vOO7qA5F+3qRrfGNKq+w11bauhY
lOkleo09l5RSNueXZJjSFoHwJxowy3re7AgTt9fFTPJGgw7nKgcIt6zSiXaipN9F
kqNd4sISFp1CT7DPvdciGewPuSFyJIWyPeZ8dUTL2DlGLF/ttzz+pSN+wkOt9Z0c
N4L51Ccpr8jgNNEuniid/kG6ICLRhdNr6SgkppTnbTHtsbkQu3NROR3/FHwb/rxW
Q6NIt7ABorNY3/aqxXzWd+UbVd49jzqs1mf34FBk0NVtVi73ElAIiLvixH+bSlHl
SW4M0Aya3eAH+qYR0bWTDPx1vHOeD42WKahkLN9VHzftTZcTrSjrRUTa/n+YthJS
hd58DZA0J7PFXTjNY0QPc0ndWVtWtiNpIadPTXt5q3bjUvQene3p1DwyFtLFNmPD
buikQOLB+94tLmyrGAgx4oHGW7M2kPehZie2VuiFI2asd6a5EcXF2UI6jx35w+dq
K0PH24AbMoTZozuHzd7KDjzuFiMHALN4yjbS6KHHMxNX+HGApZjT1OhWQHBgc8O3
s971PDMwsSUTatpnQlPd3isul2imYwu0h7GwYpgn9gNDqEjWG5rTw9VNXNTAC5GF
wfrD2+t+HyrjA4IgVXf3e42Eg6SJ1ltwu8sF6Bleh+UmMqXuyH4K/kPU69ovD7PY
pLUSUNEde0be6mm9lB4wNjBce6WaY5KtJZ16uLIMTqwUkUrbJohI1oAbZxkyubgU
VoewQR4DDvoiv0BMH6giRcry02oO/REHcbvwYXhd9C228b5p8e7M6BUaoMPUy5r1
+tH4ahOLLL8U64YqmxMcBuIouXIb8ICkERYH8OcBCTal5ygWYLtyVxFgaS+XbWCV
9SSHxtLBmohCShSTL7pdqfh2X6sNqQsoE2CfKHrC052Y9/OkVqZZGVNRvh+LHQR+
yvfAJQrOJAzQPlR31DX1ZYBgZFmtRm+rNuHgxeiKeaZmdT/07Msvgou2ep5XBNEr
vfQhObUkgOKv7BK6crfgzWVf4YSsRj23S19nEztHPNi2Ed6162gNSf1ATUganCH/
SCvmA/iB29i/sTvPmHGdM138FxFxgoLryTMuOYNKiA1wii5i4o20wTdTEY24z3fE
+tl1jaHLhNiyV6plu33NYHAxNr/HAE8k5pnOJ4nkfUcYhJNDUV13iWDgwyffLTiY
xjeMMs4nGRf22bv0X4Zl3vG0rikQ8leYeODcenDqQE9CGGDqx3C9NJDpikSGloL7
mxfIVgzmH8tKiS78Vlcx79P4+yIulgXC9hDPlnHPHQzll/t6LVrBP2Cby1tiS/k3
IifvW7be8J58YdPXi1i5vtsLZNCrFannMbFd932+sSOlLhY5Q4a5AoWQFgmSa7Vw
9/VX+SxGI4GW1nAPvDoZeRqB71raAhglRyVmOD5OWSl4qXk8hJCDogybEgm2TS85
YUkq4fRGEDvZ78a7V4lTgeZbMQNW0x6g7Lmf6bIzoxkyj3HSSyQeuKJlJZVSGfLl
wppLuIlA2J9yOvNGIW8dO3yqkIZR7aeiW1OmNrwov3iJF+/RgMt3K8v8uhtZPMD6
6kBkdZvrc0S+WZeB2KCPGRJagY/fJAylw/VXcZpsC+dKinSuhXpgBxJE8qqsQRCX
DNkvkU3flmuQO5Itb0Lq4qFxX7+VikVrlSiSF8IQe7Wz5TCUsVpWv6d3K/+94A0u
aI0Us/U/objSNLOxG42PqjvBqztRiN3xJepChiDWQSk6x59vlMzPtuXpZnp262Iw
f8ID5gNgjYFS0R3Zqtkc2+LAc/DiHQyRBXEIgwK+Ev6a930VLpn9iqEVDbCgUbmQ
SCtxowp4ucA8vhDlH1ReQunIjOtUpU6f4P5jFKA0fAODHmu45dEIpglqE0l9rBmY
3LtZ5jsVMNd9ryxBzU5aCWyRPjGsWz5Zpdd6xn4imQ/BXJSvQLdw+aDSqJ79yb5+
AjNsXh+n2FX9LhBBBqxrKrkEpJgcoOO9KbUMn66Q0O0Ho4+CXOYWVvNWc4rEW0Ol
RdaZbhZlXSrbA2+gEpriRW+02/4Tfy5xgOy317bza2f9wKl+UeBQB/8nifEjafuG
ffqjU0DKU/qDLHrZrfjm0iglI/FbuHD+Z/Aj5w/g+kee3pCGLhP3+oY6lT4W0DzN
yq1CZMqK0Q4DAlY0V7eUcsPlxazfEHjWrTkTd189qTUyg2BZmJYl+vijHJK1Dcnf
6FX8fTr0TKiPohvkxX3dLWibC0HyrkX+XOTO3LkSyX5Sk5RieqcyZTgzFEBGwscE
tHio8YMJTcTSf/r1hTb8nfR9EbzaNs5dSykx4PwJGyeRtfMbJ0dO44UIB28sqFGi
ErednIpVqNJqGfc60hbVl8DmIHdu5Jq2v/IMjw4WCO0U+RxAMR5lLsYsZAOdCGgv
Rz6DeYzFjU5vBrF+oyqfWray+1uozyURIA5F12jEDPl2JT6wyesiCgJw20SUYzqv
xPNQ2vPc9Lhks/I7bmnXn7YuQvRN733Y9YoKgchd55hK9HrB6ybynoqIZrauKEwk
mIMbWpmWmFciLqsLyugbs4xuNYywYRAmXnm0bC2vsYinSgYBn/HORYMgdh4hXPpa
T4azVDjgQmC6ZGyL6Agv/S/y/0T0BYyfZqZ6se4yYBd2JPs7EXKcY74gKSzX6jeJ
pOQtPRMVmIuVMK43g+TUKzmjINqi+3jPJJ4vsTGm9phHOBn+7p+dcrLdiUmHr9oH
Sn9RcWnY20gAIPXYCzSla85Md0waCbnHmoNoPUyH6GzZCbpWZ6AtF1vmWbyOHARp
cCPZlV1kLJ1ofSO1E4tfwcViXrCac2SRuGhf1YH/FUExYH3BlKTRuAUn75OOz6eA
A74h9xnpkqRbQ3C38+/+YXgWdpmJQpNvyIZyor71gfEkNb72LpJn92uWKh8XuhsR
I7n3NlxBw6Vda+LK1YY2r8CT+sXLjdA3+GTHXudgo8aOa2VBAamrPVKGxmuVX3Wo
CStbWucEd+rqAwa77+/5fMabadGAcFKhijTDZZCuP/MuCThN/7lbdGQouD0RfUSh
uAUJqGltmoemIzWi7VZ1elJwExYB+gWrRWJajRJdHfDvDuRu1rQuTCE+c0ZVzoR/
veLBgahQHO7N8gv9ZFh+pxn3zG1OojGZNpXLHuQz7cVHfaqueL4O+sQxwqbC36q+
YVRBfxR6RP7B/jph4EP8ROG4aEi0qr+bC7DrAi5J/nsd5/0bHgZ0i4CH2guGR21f
TE6qRUsQX/7H5uDDrV/V4ZKdb3tDAEni65arpnn+eKO+lvPmA3D++yE4CBwZriIy
+H+dawqJHtTY5/OU+Ju/sup434zpBqUN7BkN5aJRGMFsv2DlRH5wqOYKNhwNM0/C
an+YOn93ugnLvCbvBZgAjaVy4GsACqQzolahdOeRKATBKGA2lsR1on/N6zl3xjZa
j4iQXoVWc65/umyGzciHMI/YQj+/RDa0upmKGTNjd/9+gpwC9uAI6gb/AM7uO1lR
BDOEb+4rr3dq1VCuqlqCSV8gGlSN36mU4BgiVJ+vDyHmR6OX44hWt1CZZ5Xd0Psx
Ie0ejPl/ukOKTX080iztHkhX6OY5FY29j8uUIbWKUhKb3K/qc0w+PbcnYsHZWFTd
fXspcCO9YhgR5bsrG9nei2RX5eU53g8vnV2wXZbeC16SgvNkW0mNPS4TSA6P13ET
Sp+9OHxtXGiP/2JW7/QN4FwiRi+Fbp4ad54G31AORctU653Zv4JcgUSWJLV/UiJb
c2x0WSmLfNfjoPe1XsT7JzZdGsqLxwwdf5QMb98/60UNvmxJeWEl31WgwK7LOChO
94PmhHMcbRIQsRjoClAKjZtzCI8D9g9FqfNPJ5D/TBwMRIjO56vfcL2xiMl2MRr8
hUdbI00C1FzkgRdfSzmsF09XcnEpMadS0jEwftxZVJY+76Y21QvbdUsboZntvhPO
uU3Jd5mLo/eXclJ6PTSjIN7MZlKsvYSejxS1S2SDxSbKzoCxNIsHO1QJHIiFIgek
O3OpiCIQrN6ejLsQByCJKPyvoa5ybIk4PHkHkhv4uLdMGG40odu27dLxYkny43Ep
EEpCRyTGxcVTCF4JGIBDrNcECEhYNfsCD6Nc8nRKqO9M4dRg9NiskKF8sNg+cgLC
5vXxb3ydJaptAYwU055XbhBYFRsF7CXvmK9g6lNaDRWb/O3wqxeEK4Khx9jVn+di
VQ2s20btX81mSED+5Ic2lqhiPyFOSZhRwR2ji9/mmLla1ShnuVw5yQNmnA9+ggR9
0Q18U2rzZOU8nc2K3kUXczWAOIKVQ0e5a2lTKwQXwLQUbbmnX/v3G6TtwKtEMz0s
nkSJZ2gCu6DS6Mv74xM3tY+BhXl7wvz5TmgLiWABfsIXnabUv34+OacQ08N0lakm
y62FXgxsCRM13S6zw9FEhlbJZswLfQK3LJskgffARpQyaLypJXzzTjISm8BZxHmq
i5C9vkYwK5T8iwCOajXuQoxbs0DJ18mr+3R9kAvdCiCcTKo9JY63BchohPfwvAOL
+DwQ1ml7TOBJ402Dv/Z7f0WJ0jDhj7hhXEwxSAUEdI+Y4QEsEHpH6NvaZ7n4ywk3
xa7f9aRCTfeobfwg9v5Kn7JOtGUfJ6crqAtc0IsRwUz+uvUeIXeiN6yiQoUNv2Hl
D9hd1/BzDO8Du5H1kSOTzGH7OUmfWFikna/H9ZK+ktmHjIgHwYfM/jvZFKmToPaT
rds3jvtLA2avdWEsYoKc9oHyR8oCrogfOVsKH+Rc45qt2wykElQtUiWsT7Heo2k6
6nuwm5dZNKQziHrjT8RE1fBIMaQcoJQGkBiuFJgiXrO9oJB+KkxhOzpEwoN75A3K
KBKEy5ppw0Ut+GTZMrJN9QFJoGz69rCLy9g2r1kZ9xqFw3BJ6WOrrYUnkbh5/8iN
cZ4saWEufynmGFq6O8SyiefFBPIUsGj/W4vyVecXjLBiL59+7LiBhpEo+xcwsKbp
ShFpDnRwJW8dnDzyhd2/1fdKY7IUwaMON7ms0NuoSG/LlnXOrjDy/vFtZjf5tm4n
DtVPMngcadfke9JogY4SiJsOfVWFPRSuU03OTktHqsrhS2iOMak8FXzJMAriV9/G
1ALprfXb6XjXOHBKO7O36LQgQxp66ST/gEM/wUVyEQtylgNfUHkh3aWbXhfEJdpu
JVgb3k88QA+4q+ZogEqR9Dtv2SofzPe2CHe+ROvi2ILlrsLDyEBumXKXz92fpNg6
2y8jZOsMJNjcZszpy/Ji343bCQydwgnfvv1bxkj4DsmeHTHYG4Brn/BVgJTaOAVN
eN+pTjneqxTbALFqTslpAL/fzxTR3WpjtbiuaScK6Dy4LmUL8Lln/nfsJH2L52Nq
El+grz6cDyvgwtPb3ePB8U1vziLqHtjutHiB+XQODNvpjPmsTAa2IiXww542wu3T
WBqva0bPDy/OCmmNwF9sVKvUiA/QbeyfOe55KL/+2G7KPWVzhMzf/aoffYIzwLrF
aAUBk+xhj9OyoVjDMvTHMsI3Hwrioq9aMY0u8BTRw0hyUa1XDU5+v7HgNnRPtGDg
hIax/RJVo0mUMoUG8D2Z5kagWkoc5cCGWCa3VK5cxT6UZBoBl5m8wPizClvWZeIx
XUcQQ34dNRJo7FQfdGzbcAXQONqwJniKGqLYowp5blfL9qYeOn0qrqbQ4fJL2J45
hvziYhs7TIvCml7ZYYuTbDUy/h+0jQrxflUvTvyboL5e/ov04BsWIUAW7tFMeb6H
ZgZTJ+9XtAwj5QQXmNBsfku+BKvNSGYiM2Rfp2CorUV2qqhcjXgYveSAvpqLCmfI
iqRbCxlHPOVWZSzbUnkEJhSG1P4Gmnj/KZtGW1z6IyWlO0ga0sQ4TF/e8bXAalMG
VJiaGR+ZLxjNM8ck/1sKwP7lWZwRvWs/QGhLJBkxtfYi7AR/J9mV2kwURBeA9PWd
+oqRFatw+7WnMBC3SFs6Yrrj1DaFzL8fqUyuI6PN5IcKJIS0FZvKglhxODwcd7/A
whqzVf+H7icRDmpMgJqgBvBFWcX2nvmCmAFq2IFvVHgRDWcUnY15AEqtT1alLLOF
vQnmpY0VLYgaNqFEdl/FDyGUULN7q+4RA60kXc4dIMMxwJW577HGhBLxvVoRSOE1
ej7gJRmGba0cOmAOgNg50HdXdfGX5yUrSlgFSD01vss/wooJnU0cnfYXyluu7UlU
Auc9D8hlIXF6GdDP8moB65bmGjO51vxAT204WKrRLYCR7nRYthB4ck+Tv8DpiLVR
oQ5aPCHjMfpNGOMX1HGLVgkOMkxiDnVUA26TuZmIDSssQfaPvVc+/0gu89WpNqRw
351RBhFXbLfjpIHJT6rVWz6OYDFgeWdduOhuhph5Ssno8SOGS1wCppJEtO+i3vmm
WZg8um6rbBbSbAmEhUozERccPGy0g++2C05YSmQM6iYC66Jnqk/AZuiSjnMQAgDy
bPApYehQj1t6mTzL/F4OhFmq2qpWwtkctXuvYOJHtnjSpI0MlTKgHckcew4R/pSX
slfhGDPLTvkqLU1ILhNhGb4OU1+L7PLqDqSZYx4gVU0hG0bI1JR3UlyoIb9cOzLG
3oBd9z/r+IgNpMtIi3NQ7ATMJnKs48SZ9924McwX/Je0KJZe0REABYiqr1XR8Grl
h4MF73qYxid+V+pia/6d90NDJGWnQ5T3HNc054Z16i095kZm2N8jOEbWeSK/EZye
gIwqwdUQ+U0K6vTdDSQ0B0ogpnTpU0jXPVp7gi6Jdn/GvmLbox7KrbKu9T7znxL8
5ro1pbqxVfMpG4VttDlZM5Xwi7SoFCzlkRlMhz1bIDcgPYgt4PKlrWelkwhMmXs4
npigPH3ZAQHfu+UGKqnIhwZY/x3ZmOfhxsvSNuzG8AShKpqcWpkMfuVFY4wnYKbh
q6cZUSbeYz2GJlxGzFdAFBvisnHNTrpvlSHPT8iwt5tO+CFpTBtaU8E8mxBzHNuu
OO/jkY20V8DbW9ru/psINFKx97MYFuSxIBqVMEL9tB7iqNag+TxWuvaDFbMnBUqY
A2DjLmKCJhoNA8sydn6VD0AGq05m8fnaMgY/Kzp666II9UmyjM7Y4yTJTZbfWGAd
Q9z7bOhEQxpc35ar2f9WhYSinlt9DA20lakLcjX9fSUQjque1ssHIBz3oBFB+OcQ
39oYReAXUnbUih2sW4E8v10iJjlef3k5Ih5/QQFYusABAxRaqeWCOgJ+e1lNtLP5
8EWvkaUTS4wn4/IQZv7NDdTKbKwQqj8AqORIEZn+hZqEsu/gJHqkNh+sqtGweMbY
D4gVSQgmVzD1Jjz2+MA//ErG1UvmfqA/A3D8Q4dQX74gGoLKRQif2mS1DIVxXnQh
orxRmw7+GUYVWOg3EdyILLzf4DrEmZ0JLqZxWL9wrh5sQ/GHwg8rmONuhc94rEI+
BYuO7gSV47mjQ6v8pR+xaJSIIc6IOJ5wgM9qZVfy4DH3a/qEh24sKjuE56ulPpHR
kFlUmYdhWaIA8kCPAvoOzS/z2QQa6oZ1Yft6psa3hUr+sAMTb3zMkjoqbi++hVhF
Ox8f3qUmfGqUwRJsR/CSwQMeXOd9iMdfzPgZwPUlDuZc9Wes9fWaCkM5sM4OjCmp
990wl2OJ+64Y3qcRN1XCuak61t8TQD8ptKixmKQzZgHSfgc5QdcBS3kogtgMzPNX
1+qucU69Bm7O1DVde6v2Rj1qAE0TXNs1B2fHnw8qxGcUHEnkmoWhJ1Y4dqmq7KRG
FiPp9bVKUx4X1HGWg9/dOO49ft4x00JCOAfXtZ0XxEaN1iqYkSX4hQhlU7+HfEHw
cOs6qmTodJal2LYXWVO4aPbR+Ifb6RJrep2y8Y30C98ClRiCPi5EcPS6ZEyPc3L/
Wti1vFbmNU4GWcB+Nao9IKHKicXitUQoWHf5c7Hjb3ffNBs/bHcIEfIERPdCYcmR
UBXtnsJL90BhUAYC7FO6HwC3R79u9WwiSb/YRD5KEa9dPItufGd39lMpDF3zd7jB
PNHHW2VaTTH4pe1ruNG2TAbQAdp59pbXy2Q+mEJrZNUhNeIdCUX1FkFNNm8xyJYH
fbJAdz8eeuzXk9vI1KkJDR5IhV9jyhERbPx41VtXsZt+u/vxNlaDL20+WOdcmWeI
D65/3qDQyivM+Lch17pbUGR5WKb98HPsGV2w090kCxIohSleiOW2eMJOz+bswTli
aE1q36tApRfwHsEnovh7+XkR1mIp3PUjq0AjNTAaV2hs4QbFfYsM8o7hG0HlwYWy
4qPVeGWTCFFVifGWM7S2CB5cHoJqvhHFdcWfoCc34iyF8oN0w5QIt6Jh0YQ1P6/V
5MSxhtRUQHePTICZxTrOATGOi3jmHIRammUbNrtRy5qxwaXtxKUq+z8L6FdaoOV9
RcKljZ9/Wi/osldJJiOP+GbAbDMkvNa5MVZqCXxr2NPcMRcnMqQT8T47DwxeWScl
nSzKIhPBnU978cA17VymqYag2IA+hiwKh7FLLXkbppHfHES1hT4gtFBUmeTrmPQF
3w+CAsD8scbMD1P7XqemHpObosULAT2+5+DYP2fNKg5lITyM1jWWSn2lVMNphlIP
Xv2NUxqWNLUZFQ4rNR2G+80fVrR9TV8NsKVuTEow27SGnD17PTZUiuhlG3ngU4vl
GH1BhLBx8zLjIu3fltiEcgKA96wP/p2Dwi/S4nkDnVmAQ0FjFSZY3kAgrmNt/Z1Y
TKgGUmoE45k1QsN5xB84nVWDwy54W7rN4HM8cBcHhAdaBP2qGFTKNaSGEmE6gmbc
YLjQfE4IEVRqnpKz2u780fDZ3U3Dfw1w0xEowOboobPk4MGjkA2u/8ieZlRb0zpb
4tv7tIPH+Q8kG6aNuEjjAZHzr/HZvTL8y9lyMqw4r3qTWGp9ZQI5tFwo5rwfgetj
6GM0K+maZgY7Ef++IYXEOcXkIfLIc3UZfyOCdgQL5/KUeG9M/qBSQytn7yrGcHKV
WRuQ3ZIMgACX6kbhzQZg2qorRVQlWGhElsqz4HYPq3xi8koyXX58UToGin0M9cQU
RhndAq1Kjjn2IWrrRFogAWlh99P0mKPN3GEx5cTYep9avIejVogG7ZowDknTxLN7
0vH0jcNOkAc8fYcpRCg4JGN0q6F0FPJpynYhIzz4z/Ja10VzwbEaXYpBTNv8VIJL
ZiOFYvn6/FyEKCiBxbNhqIp/S2NU3ZOhcQ/hhiu/QzfbEJV8fCxwslfUW8NIpWws
Cyi1cwINxV4mENUFAvwyneIXdS2B0jdb7WrKOizfECXl4hEggFHBww7qt3W1pmI3
cLiEClOXJtQeJGHgqfK/Z0efr6QGTcc/XfWYKuqW35ZbteozGDSxysvQZnJ4DUUq
DfeHkjRA29mxOYk6t3h7OdYwdFtcKof0WNr4IJk0sXprlVOKl02qHkhXQcyQvmP7
kIScCvu9/1vVGhyCxUMPaHAzCIW854dqvy4e3/1lMNVK5Mz/b6c0as16DVdFzjBQ
bTHsNB/EzlcfnH6hItQ+E313UnJCMCCgYXVU28k0KWrqJ+PGVFkowSweTuCfqD6G
Z3773FFSODQcVN3MUBWDWneKIl+EsDK6hFSZqkfUS2TUyvc10/LMcSXtmnt3y7iv
d0SmiOV0I+chiy35TcX4XMj+MxRPTowO1TAac0awYzFL7EoIqPPZFML4x7Aa71Fq
iFSyiODkHHUseV1WvZ3tSM6RBOcecrDioUmfmKVryvhCC0IbAxvJ9DWAn1ZPb7tG
hxiuHKeLXh7OQzBkstozLuSXxUJJGS+/Yt7W13PpqyB4r8jUL32peidpK3+R833c
Q+KABLKFckzmIdJyWSzbzWPSy3TIptHPEKO/JdNjx48FvPYioC1Gth4g356IQSW9
cIouCdKv1AdZcGN5tsu9tWUdMTF6du5it1EinQjbD0oRUPQJjjRphAfkb+EsOZBj
Qh3b+g/96/c64k4Ltz6e19cggg5EKQK67sdvGeNI+S3B+8cEzz+AxKccFyVgwbLn
irlVIDXLaBd4/wZtjkVZtz5YhwMzzOqrHWda0Zrtr/XShU09nUecaTKBxjwkzVPG
VgyB9oKpvxGBkQaEcIj0uM0nqOUe1mzkIn/OQHa13pLEnumQW9OHR7c0WN79sZN2
x3nqiIX5MEzjfbFs4NraAZ7c8ssrEV84b9s+FoXxcu26FaPAvvY59B2j9pXICS0M
sNsn+gt27DB/1Opby8n2NdTrycOMEqwgCwo9jsm8wq+NimvbhAVRVRQ0iEt6shiJ
LDm0hKZcqUG6LYXlE8JgWaZOQQN6ZH8CCCk2gpeZiSWInZekc1HITn24L2ri0HrJ
7/wel/Snuk4kVVVS6Zrw1ltO3u6zHKzIr2DdfHYjrcRvz+Hx3XXmMpNGWr+921xD
RvZh5Xj71UfShTTzXBZ92bIpXcsCold3JOo+od9XH4UTkewuPNTXO/QBBq4ZJyH1
bXhhgQGfmMeFsbpqq5Lr/eXfbw6aiVE825fPdO8S/g5NPgPCcFYIVDDtZF8MuOMC
thlluj+gAOqL33SsSzJs6lPaJFKnzbxYz8QYAbANxfM5W+sMB+wQTJ52DdUDSva/
SXwYKSo6wqNtpvYzH62mKLuZVOM8YVfW3g8IkUjliywUHidgSSCQeqKe5tKZgUD0
LO4tUzBMhrJndexgB9IynQ18b+iXsH9ZB+YZeJZxuqq8wGAV3GqNynUOo8WRYJBw
32bjHlJTCU09lD9ovr5qqAcwB56sYNDzFl5+lZW4ktuo9BeTVj0z+MNBzS3Sne4q
UraWeEgbiOzuJZC+SIl8llc8O826SrRUnymBcz1e15Mv3ZxiXD3Hz4LKv1hD2t1T
yKsDhc1uTcx8U4CzR+5XYfCbRrD4GDU4T30rqeeevqxE8skcHTc14XsqaIxco6dh
GlU2vdN1DWlZRkwCi7Yl/ZAfyglU72mdyRAjuxuEov/NAewrwIFWO93cXXaBhGXA
NK77kTpnOnT8FZNmK0NbQfQ8f/VTMwsVDflAmdPn0EITPr7nTIYTgAAWB5KTk8Ub
eXEIx+n0EhzIZpXxd6Ghtra2gm7NC49xGGkO5kJFyCE7/C+WJ1yBdG43P+E1IQw7
uB1FdsuIuEev0QLt+Qy5F6vsM45896vbq9QXkhxOcqlnZTNe8zvKA0jwlIDdhNQ/
RItFDpzsHdjLPDj1UB9izm/M6SqcQ5IYd0vErWDc30E0rkrTVqXcV8vOHYJMS3UM
5/TZ5HLHH2VDqPnVrqxZBxrMgz2fCAwladR7feDVhu8XTdkqToGWtVg1xtaSJTL0
D9TrPKtqpSWfNWLNSz1qRxroO6I0hmJQUbikx/ifUkedWd04LgA1tEG6LetqhZ+G
SFE6y+fC1+19wtZ7+M9XgIeD0DpY52OQv/Pnq/0+neHilTBHhbEARisf678kpBCo
nTb5wKrLdeJi5xn02qH4OMb07dP/+ctQqbmlNWuNarIKVn7bNBDaT1ErOaov9G2G
8ItrnZSb8CXJQS9KqSHkRHygh5zFeCcGt71nyEHtuZw7bCALGWhhFqCRmjSeJMhB
ZB+kMwAkKsId3VS5klQEgOnWF9BloJX19BBWFw9L+2A0bydaHW3aQaMBnwZm5eJb
2i61fUmPGqbrwwA6IckczLfz2QQrGVCAgteq0mYMjBUij1OZ/9RO2PraM/WJIYH/
EDnbieHGMssOqH01EUot5sj2P5DqiKsFmsgqigSWwBpnJMSW+PqtybRdFwTaJivG
Fdk5l8pNPfg86qWZQ+EA+zU3YA9BBrHTbHQ/DszMnbba9ddtTKp6Uyq6s0/K1iAt
WtaMn230xiMIT8x5G9tPIfJsytQTZGz0lKr48NymuoEwHkjLZ+Y1w4ctYKVEihPd
Vx12UphuvXfrb0J2gbI8y0HOXFZTlP5tx9XJBHbeojaagDBjpYL72lMCOEvk7vgt
OG2ACgiOrmQfd1AFX8iSMJsInvz1f2Us4+jr46V3U/nnBAPILQYlnNI21VuNvDaT
leKbwh3SZpx28Zn2Q5JZ3WCjC299K2gCEefI9XLXX2+y5zFUxaZsJq35Tg7hdnqA
zevN+VQ3bZOgN4D5CyYsh+Tk2pmkJV368qF/JA5X5HWuFduRDxBYTjlHPfqEzigy
Mqdy4pjt92Ya0pnQ8lA9yVDaR7Ee13nruPB6o8vOe7ngxbu5ltTWV3MQMBDdzeaw
zYsbVmX/dK0khGp+MUuaeAcc8RNtDBY6+93Y3QhyRQULmDLzsF3K51iKK/CglS0F
lFhzjCIDlKExDLYqPV8Am8etqtvgR1zgl6U6OkgV3pLfve018V3l+0tm7xzo5vtl
kzZOSBM1ZZrIOrfBOJC17SbA4gXGsZEEKUQKBFcwnPY6jZjBYiAjvLynBPPE6wi0
W1K8f9WjFhz7deGGPOmj96WhiIOR4CZBgJq7U93LaRclUhO2mOUx5LRFLxQ2HBLO
vAb4DrdnDw5nTL8N88PYui7Kq5W58n+KzYeuYTffBprBS6xVrCSsGdJYk5uP29ju
49v6DDnCCzqI1r82RIIRlED2WrWKDChNvStDjmhlcaqct4zzacqym0hPaGcEf7ai
EjwlmH12fRdbLQr6S7XTSrD7stAz8ionxzEMJab5pPZ40G7U9pVSfzg5n8OjBw4M
JjO34J3h2ZQiY3RdIBPCxqZ0+6ZAFzp+8dZ+N0dANgkC+vnwUxIRziOyziGPwaui
/0CeOD7FXg3/8Ek4z+b+5hasHhOUCXtJ5xBrRr9lM9Mck/GvW4AxjKgHWp7DHWGR
/QZCL83aKlRUjsyKdt3VQpidlKb1XSLigtMgTHlcUucw4ZSAKgS+VgcovI31XAKk
T2bbx1YQ7A5dpwILq9YQEqaZLYPWojIGgKISsjA+o7jaizrVcm3g9Cd4FtxMQ1WY
YLu5R411ehe2+kTtPAEl739qtOkdKdevjx9GL5su4XByheI1DixUaCBPvHWBQ74j
EC+cL0kyV99FJlvc/Qd9vIU5ujB+1jjaO8m/eoedNdI5uMWr/Tbqyk0cRzYa7WjZ
BB58LpjnsRHRMi7/BEutPeYEgbYrhKyiY0/Bbu4aFDz6Wa0t8nW9Lj7pRmc3US2T
FrWk42psu9tqqDTNE0zEIVxVZC9qluMu2Zyxdju+lY0kchL2Ljmht2hr21hGM5WK
UbFszyYYJ5Qf9OkPuuLt1TE8acUE/0Jy06Bfif2tfxDnF7WhIcDGw2zn/6dtQI6D
7kPYuAwRmCseE8OK14C9keDkMg+mzqiEqp75vJO6D0bnjUrhE4440Ss1laC4U3k8
2j7CdY7fQXcV+VKbuSiPj4gJE3r1pPnpLTMIW7kubY2lLioI9FMWTX+g8OMh4m2M
ac8ANiq7nuslqCiJBqvdlWEv5Rq8g6t9IJBN8SKbaZRbu/OUg0xMg7k9iv8YU9Tc
veZO+9kCwvW1P4hy6ftI0xQtyvvuRAyW7xE5CzFz1ie3fyJN0xzsZDdsQlA4t/CK
lRIAc0uUnJwpDr2sSLIbmPZJNZY4cKppFRVUWGPKp9yoWuq23xyJwXn9bKTxBBO0
0m/jeBRmn8CGnjRSOyw729IeQwAhRTHRzIjK1upqmHGfyoVPJ6lVWB5OaO99yfxX
vIYhpzt8JXgyxWIcV2B/U0A4t1ZQNVB7DrKxSJLs3z8/HA9MsBt04/A3uQ4KD36s
GDTdXWasSleAEqMirpFpo4+LyRJ4o1bSyYEtXtEQDCjHfGI6zyIL/n6ilrHJjnRo
W25n3KJkJwWheO9mYF0m93tGJGX5UVD2tMrO6hYiu+TFtzfhYWQtPWBK5Kob/1dp
oRX9hwOGLRiAqx2GFk0106llVhomGWMsBzX//6b3An5ZCoGOYsf1zdJec/E1JKOn
kDozuVX2pJOkmZLRnRNOzkgt+EIA8HAodMiHV3bjKfDKpm72R4YpH6x5MQu3aYqI
T6ax8AHpdIUAkoZfiYGC3T8CLlHaYt+//IzSqzizx0lIhY0WA6ZNzeSir5vy6XVw
9IsiG40O62DPfqOy8d0Tgunoz43bThAy87saFisW5E1ziTolxYcgUkO/i7MKpBOz
xyTZdx1c6Q/0Zd7+mcWTombDycFRhERHBgsASRKcS8tEkWY73grEoo8UHuFp77GC
hN8TFT/FTGWdJ1T/FzWvWI4MPZudiRKcnm+W0dphuRnlS5Ezwq5ScILuY2U6O+XD
Mhepu/8Pe9JTzIkLr9C8SheMYdaweytRKFDH27hqeZLAHK7h2QXgUwHMrvJINxry
cl9GjCmJOKpYuH47ypTyVcpNZj2nbTxLP3aDnfgh9GHjjvrUkzffadKLAwrVvNaZ
wQy/gfJMzpIIZH3uSLg3PUxMlqIjHMr8HD/bYonU/09RhHh/dmNKqTxB346/zw/z
jjXcik4ZWvTruiUI/+rS5OYDEdW2Zv/GQh7qYhfiVOPD798MEKCsx8PHMDOiTlAK
Hpt+8KqJ2pEiApH00x7FvTSCRugDqzhkId0BJrBXWCN/dRdBqdSy1mvDcK/uJYcE
Ic4jOmDrEsSLE9/HUZAdEPMXVxWlB2rQAUxNSjZVskqHOcCffFm58yWxDpxbtVj/
JqcvkNtQbdNk+L6tYVVxoNWrjEaIpx++bgnb1peHv+5+2Xv87pg2GHV1FG1Z6lBh
p+NUlA2ZQlUqu82E0X7lQTy8tXaE3kt66HsJhgZRaBCJXF77+OBqjn3rJ3MOSyvA
Sd8H7yEhpqvWGuc2yh08UlwR3mQN5Ju0Y7A+D+eJwR+UKNRSvVv3uDG1x7//6O8t
m+BzfmF5lsmRes5TfGx5mw3icVG9InahHhz7bZhDcnX83P43Ttu5OnzzHK4o1M6a
TW2lDx8ac3afDkffx9WwtMkjK3aSQHjcnnszxzzDTK0upqLz2Oet+DbHj3ShnhH2
5MUYhaFgwqof1VhDTPjBo2ySyoz1AuKYlt3mv/b8lenJOz4VFErvvpKysuyKR6UF
8S025iO95lmyxpkxWQ95/0Sp9k/XLnkQhswKmPv1dinJ9Dw/sPul23zG/Ylrh+bm
9I/QJbICGyV0X792rt8siaFCDmKkR5UMTkOogrGVdV4bm+xtNXotBXmY2GoGqfp4
AQP1xm1CxRW9wXkUEsKYMMyg3qjj7EKQu6Os8NMedGxMNOKvZ4LciDRqlFMLWSKe
wRavIFHtbjTjJ9PDycK+GtFgxcWR7E20s3b0gqObF63nxZtzUp97+ujyDmh+EtSZ
zQkFDAg4OgL0ihVuwmkasbyFWdy8wSspgmczKMXR2YpkNS5Q+LvH1hFPineSAIk4
pfLJzyCLlmaP03i80sWOe4wrd6q8vIY74JvVsFMLFkMrMoDDARpvWAYIWpTw/Pjk
rzD+qDm3ZMEcFanKbt6fn+U95PFrq3j5qWNbUkfg2ByUp0XGUX+hzXLynl0WLe7S
12GM0SS6PBW3yJJRaixWzWRlYHgV8CNLGgdI0IBNxWd5mPcMevpgBPW5ftdTWF56
L+vRyf1k5KM0FT9L8dMqO79S5y9JVKpBUp74YAD32Yrifu5HL3fu25BsLMs484XF
KUCfSOnCwlq1U4S4OdcHRxAHPGbyYzSru8rCP2outD03vUtp4EQ83izWk0AvuN9w
NsWqvDFSBjRGxLcHppo0x2cKVmc1SxoBUZfHCXy0LYK30bJ2+EwlQ7Cs5OjlyL1L
CGgL9qRLM9ktFJxkLkRlB2pI14ZZFTxlExIQXNDnNOikE7yaqOemWsa+H7pdhxNT
LNBZMO0RQ1Up/e/jIMchLZLztGsNyoMAfFy5NRFGKX9aCaHPUi9UBpinfNBU88sp
Qlgd2o8t+fS9/C629zZMoufaTrDj+hDUEF0BX+jSqi+sB2lZNovGpiiVjfUWVRd0
xYbBtPmMV4IPN7dBxGVRO/2mtzaZooTb0jCoTsQPxj9Cn8Ke599vAsN7uUTFwRXu
nlIcnrJKCBWe58kj9vcG0AatbugdsFAWlJzhQHItdc4u0biatJb40K+t+lrd5LF0
cgXZkh6jVr6ONv08b4BN8o9jux2nZzPUrwEkIiUIjoOeLGbzZVC/0VmxKFeNHn7x
mOazobQC/VAVW5Mr2Xfk33PTtcCWi4Rb+K0bS5nEKcX01ZjkcKfBMcoifg4zBtDJ
Ci9dFBdGnHPx57poRhBkFo4gMXc2aHrlCObodA472JoPsEO5vGy++Bpdx1Nny7tc
kk2rLs81xF5VnIxrdnYZPLZbrY6xzQwv4dfbFcpC8knOIhJGRIYMb1jIaZ4E1ZEB
fB24SXDCb2Dh2xRxknT+ebbVuUWOalRG3spJwy1ZLSRZAJnYWJ371geCGA9cHABA
CXooRMbzP1pPCKDzsp/C9c2RLFk0nUhPKfN/ciPgUu3oIVwTv39khzy1jDgqZHL9
kL0YZExUYhLCzQiu0sWRSvaQ4VPrC93a9GyED3b2WfyPQclH5rv2S3WcPOK7BoKX
BuZME0+GcL2AXyuMaxU7wQnkBRH8XfUrQ6A+Sq4n8bGSU181+gr8XmlBfUR6wY/Z
vUqAYKQrVvVRqWNFygOGkeAlCPhPpLNq89FA/pCbj0C1j/eCMO3MFR70pdJNslCo
E6LDNyV5TQAALCZDWLlfg1bMYKiGuxejpGB/p/lcZ0aTzTmLW6DItjWNzv2JvJYa
oafxfRI9TMXYBRFQME4ZtWBBUYdCkjG7tpB4jDmSAA71e2t3AyEjiQnGOKvRTSh7
1h9QDALVauawRU6u+LR9h2mH68aN1haT3qGgynM8l31TJaKqeyrkIFPxepiX7mbU
P34QWIqrsXMfm4YZ+Y79K30BCLyPg1Ku9PcyGE8JjhkSxGKb1y2GhMN/r/1D187/
GgEksKohn2UHNap21XnC2leU7CL8u9FtZ+DOJ52zvFVfsAzrFoa15oLOk0DUOrKI
PLHlxRuK4U3Iyxh2qe76vnHaer/brDDOUjECowq4SykLNnzYns84j4WB0iOjC5tN
QY5N1R6doI6xr6bSB6NNNCHGB9xWZVT4915sltv6r8JgG/b0hHqU6K+beiL2qIrY
bMo5RKnVHfOsPVpZKPglGoozAX81Iqt5O0MWtFZFwXr0w+tJPVPT0DuIvgzKHLt8
1Ju7SJ35Hr0MARL7xNL/bVka9osmpHERGzAX2QdYVlEC1Vd7PmgShOApGGJ9PAjr
OcAxOO5R7H571ybnvgBwTZC5ghAL5OXo2mZuSoAfM5Plm9mNxbgKXm6BilCRcJwh
g38yb40J5njvlXOUjSD+MXAKczsgyBQz1SSy5x6FGMhrpxpGmuruch0nXuOm/1qo
ZkhQTd9U8dW93mIJcANFq90rOWBX6QXcdSSGQU9qvbUp6CUyEJ/sXL7ndUeflt0w
GgyNSisOuvzgAJbA/W5298ofaYX52lOcQ9Jlrh2zJt06+ZPBsIv7CcvrjwGpySpO
S3QyBh2LypZMJUlA9ZI8ZN7PLRMclBQgGednr1+IBNgrJ2hY5PI+PpNi/RR9mJIQ
p7CQkxOoDXzo9xUzvwS6osNuTqnYOYvwlKzRMEv0rGUEaGJDusxhtTJdIvVQfhCs
Jbj3vbSDc4QLb11FZwUiWS3oeL5+zWhy28v5LMb7x+lRmg67qljGACfzuSbdNawh
BRYoycKakW7xXhZyzigUfFqGFfd0DSsEIM4JaSaSKBZwlDHV77aA8FAl9SaYs05N
I5Dv+qhpczv5U8okV7JSq7SN4ArpK/Ee/h7p3I6iaWtaYoJwEdWV+yjgKNnTToO0
3mzZCbCG050HD7gToiMb0Ko0cx3yHfpcZu/JDAni/yKHMRuRB/eputq1T3thWDqI
zYYPW8n/99lhdYOlm0N7oDayRwd7JeSRgS3tgLUprL8rZLJg/qw8NgxROQztibdL
pLT7yHWyaTNii1rRsTeNbAm5XnOihgkx9tU5AHSdevuipI415n2Krt5DYlSBpKA2
sUes/jx25/T+9K0MB7WrxEMBaVx81po1F+O+5xYF81+b4dghIpQpTV093CW8BSIb
voZSVtDFSrd79RGtl3x6iWdj5UBy8+QAA4WqWXBMewjrmXo2NQ9pbclOVI7Jf4mZ
Tx+VtEg6LkmfrAvUA1qN6c3r/YFlz4dp2QZgVc1AhFKCoKi6KuUNOJw+KWydgDEe
UJLBqW+R3ppq59LptpzvSEIYWTYauwsguHJGbvQyRD3xFz6aVMPlFOc+8rPSM1jE
7wklTwd5qweVzX6qdYTWuB20CukCNXG/GbwK7OZ7M4C93rDd8SEzbd0vRWtIvs32
QdxLHR8UdKglKC3OiXiYHqInT5SBuAWmsbqMzj8Kzk+Tpmx4U/MRWe7V/fqAGo8t
az+CcCQeLfkE+kKmlBaVzh1o/2gVz4o+HbpFNG9Zsa2uV8B/zxZobFRsQB1VnbM9
b7KB7fO8Sc9xLmAC+VlQNnvNQJvPJICo34usxjc7rD594RHY1Z0K3XcBo5hEMvum
puClxNY9ZFjRQZYMw5937QigwB3tBZ5IyOZyaCA6rNJD94WW0JML2kynDtqyhTd4
XFnxtMv9Htzn7OJUhT5I5YmyRVJn+25tKxZRaWdb1FWndufG67oxb8rUrqB1FLFn
nrDwHfoHhTuPh5wZlM3Dg6XN0BeP3aRRVVsOgEZNLkCGqRkc1C+QelMBvigcr+Ag
oAaVsIvD3yRsTeVVcleM+8V7s95xlsWumlvc/DpqPNyUrj5sX8rB3mNlGn0JtvNh
p0lp8HL9mtopix6w3c9xOx1j3wSfN/aCFSQPN+zOU9Gz49luLxq88r0KgUaWPUvi
24cWgNHZ4TDkwvkSmRvKSi5mRClk/EvX3zpeCf9g8kJ6RR8kwX/4RGMUNIAj0iUT
k5M+coJhXj6HG88uAHoUonMyWn0ZBD8jnr7nVw/9B9IVFaGQuDdXTIbUMSK8busu
mW8fCpGsWqWM217iM7ZY5CJ+vLdEj/DADxd50Ptw/roW+xS5XQjrw2I88ujzzJFT
aoSxqllEtWhhGUKu0TMQxvCnigZzCcLxamgRGcW2ZL+MmEkBSIiK/L3kwUHCZr8c
7ZKlBVnuaROeTImrVq6hksU1AJmYEDSGiNfTkfqhNajFV53vPbuST2ExKYnotMza
d6Z3FrZkMkGxnQyTAUsRiVsVS3T7CYht39TPb7dote9Stl9A0j3NDVGATQ1vJI6Y
KlYj4TW4382sUmjGiSUiPlRgHrZ6EDT6ycsAoqlC26r+sE2/rPyMIjptSsxSVeKt
otCI96B12pQwQnHyBY6xzDoJW4vgvf7S2Y/s09DuJm4Ad9wVcoJG9hqzcRqkrDTU
hdgnDAZCDImIZfBObrlWVmgrrSLVbZnzBafOqeeYS70+gateSiI6PfOrCfIVVD5E
2py0r8j2ODanJjFBiK7HiXgWQu5QwHEmsPnEYyTJ9oniPT7H7X4BHmrBAHg9aA0Q
x6ezhvww2KUY9CpoQZ6RCQizNtVZ5z+hi+Ej7FaKI9bt0McxcuChmkuSlPXYN6A3
4gZf8tgTFJo75QgUwVYTWrOE+jEOdF36tX7hYZn6iiaHVB+FovJ5UFXl+MyJ/soR
XXFMKIJrTIlagx1Txr5KTSifTVJaeOBB8zZ+vwKZI6MBHspVAxYa8Nq1PW0d+HpH
HGEsfyErHVkkP7ZStA8KuwJI8Vn9eNmZ5yAkRvvmKZhCDYGzzSTi3ZDh54fPPIqO
y3F0/z+kpVA5287NiXKDhB6vcKS2RyKPvyUdRahXOgEq459oDTvVlix/byBggLT0
VXRhWh+/7R4kGvAtawk2MX2F5veymr+nYjDn0uj0dSmUaSSvl0S2qzO+dM6N1ywY
TEzDqNCcf3iQ/v0g4Dx6Y7M+jvTP9eBVs+LIoIj8mwKCf8UhXjGcxJysMEbFEDoP
hF1snF2dYGbZFbhG3clA1YQTLBT7Kt00wgZm4Gg4wuYz8hEr5/kzkSxdPOk4e+63
rUi4aPvE+9VUSPAPL2GYgdjgjxZrSGOXC/kPjb8Ofqjr0l+fSY77SjweBQNK5has
OZV7dtZ88jVaO4uXHZbg//KpG2vJxxEmjjqZ2OtJ1IGo8WMMvO/LkgU42D9MyYVB
wELtj0CyNMNZX5dbRcbX1XsAdjcj4tuVFHgUdD4pRCA5ye6tB9vWWulOO9Kr7IjR
9G434fIMk2Xq58L64Rfbv/uiQGePItTyleINqxx1onjFf1RSne5GyiEhNt8gxLto
qRxmBgq/OjxKbzC8yKuqBoYnvCZkYBVyNJuF3xTFFE0QuAuyv6iCcG7fu+tkIrPE
xpq8lfF4qsYdc7NaBgSuNoo+/3XqnQBXn985fOTOLUW+m1mCrbdVjvM4InvWLifR
BWm4fC3zrXjCYCKnGSqChLRE+J0gE5Q1PUaBWQ68Bqd8PtNiZaw8d8Zp9RB+gqF3
peoQ87HB2slcpcwd6x+ay9NMl5xpY13yruhKkmzAUyrIGceWehgHuVZQxdoSvvwZ
Go89DyHNqDpC3sAhfieE2GgPHxCO7p/d5ZO8bHR/XHV0uEhCty2tOUCoYNcJ893P
BUFpxNncaJ7n2AzBcWjiQlTc/U8kG94KIHaHPVN63xST9+c30WGUN3gXt1lHQpAi
dLyTJQ0ExHOeQA276eN6JPw5ZJmqvY2we0zdG5S04Ag1mwXQnRYDGaBFovuZM2TV
6ikAtdovnGizDhqXWt6Mv8eI6eupohCIBLoy7vfMG2KPPBR1+kxJkrvJPeiUrFXm
BSZOSxXY7KpGVphilXdSlsk22b80c67DQc0sh8sXRzubt5dbgKeFlnWoiJ5fjhhZ
DQayVdMOlUTBvaPDZ2TZTjK/MDVyimrjh2cS6FZUk0Pb+Ri5D6UWM17indz/7C7W
+XstceHzbkc0t22Eqzj/WjreVzAo7UbKqnjDxqUNsFuupoiR/fQYBqYTJL4uQeJj
oP1WB8y074XocDWs43hJjeiwZot6G0TjflquVdc4aCSiP8MfpMKPCTGR63G3O1cY
ukebhEtFseT1n4bUD63GVCixhndXMZXXi01OK+zIwuRnP5P5mWnh1ifCb6RVRDZ4
pyFQesot9HVXyX2urfvrrZzoycTF6mUAYY+mdzAi/p6VAWnaZeA6tqzLmCtG2Xvo
eEVlG337M6RTCP2SjUpQJM0NT3+tAFts7wg2l5sHcZw3kVOwhzIP6hvcgra9wbu1
AoGm0lo237gem+JYOzpS+WlJpL0up2AGB6TmEv5OcxJa0FM60tDj59BXlGQs65hn
EEn66iEuKu7PhdzOwNv70GoJbvhbqS0HkJeGNaZTlv1PPpe4D8hTNUN2nZnMoH2S
Tv2mlq8/EHL+/yi6oRULEfSwdhCWNNyCE/iZ7D8XGTT5KlDLkdmoCbFOiCuZHZY5
XaV9/e/SR5qcV6L/9CKzQTvBl5cA5P7db7NPFhDAJTy/c2QPn+Hs3IieQU3WCFjS
e//xlqXgGFoB/MTPTdPpM9Hmy61e4ORaID7+n4bXNxFXzyXESAy0b/JkbsYerZWj
NKhup9vCYAucX0HA31+Ro9Pg7Z4eHfPTgupXO0T7fM/5a3dLbn2i+RAlQY4KO8vU
T/ki75QVeggfXM95uiqryqvN4dQsXRW6wpGxf/BYt5x2iamXD3pn3doeP53vaK+L
lzgPQxFfLmst4bwCQDnopOpvBvKWqZ9RtPfDDsHXjE2+h7HOTklG0hqhhgccM7Tr
13CuOY/Oknfv/J5YpBZF3uTE7KNU5m4Zd20pv5MbnO4E2Bx5BKGK/4tD3a+zmP81
UQ6MF39jn6et1t2ycZSivpTFu9l/LaAk8fm5wTuU3mtGBhk2MEomU/A5MPfR7xIG
TWUJk8Z8ummOqMFy0uEZz3qH9uYw/VGqQqDMYKgxPTLLt0+zLnoTqWfUhmVG/M+B
n/2zvtVEL5gDkeKHF7Pn9SMMPYCET8zzlDpg8t9xZjlAjKMGJnkaCVJCJfMJ9bBt
u/G+qWNBHV4/ORCj8EJRhJNsVfZGbu0iwfjLm5KlIJ0MiE/to3hXWH3BGv3je5go
RLNgXT0/YcNJJg7FbzVSMfFk296ZnpWpZGN+Lesrv5G3VfmB8Z9nsmQ6bA3i0Q4Z
Y855D8RV0J+x4IqfnvmmzVz6PSFQXUZzBh+UxCJi/hx21WmaaH+uixKlGedVpIDH
wUs5WrWC42VR+tjsEZD8BxHtMh2XTT+6Gfqno6fMPsfa3MkLgX7/355VllShIGaO
NXm0g/N7gZDd1j9S51cCsZqhTeT2qeoGsnyfNkfu7WfxBAaHja2guWh8+eYTTPxs
GN2SMGFzcs3hJjztBRxVq19qMp2S1ffRVe3rJTeMfznc+67CcktK1RmmNN0g7Nb+
SII/gwX0/Ag01iLx3CD+fnrCPj2Qv5emjhTATJI9R2dqIlF5dY014YiuwRKqByCf
py5hhjNlPTzhSNUWZIPAw7uWaQlVnLanVddzcHquiskfEB9Q+wvX2guSqjWHGhuI
1JB0A+hL7PMU9HwOhVg1KPXO4Ite3OWNqLZrOzW+No87qCWgwsa5gRpiuwN3k5LN
hQbTh63KLRukyt392lrq9OflmyX8nZr7ecxOscQNNcMM6igwQblIcDvPcOg/douB
7LuFm8M+21xRRZ88f4lLlUti92BpxDn4myvxKqIWMuT/iuMsJll6Ei8s1tEaWXJU
uEHaW0H15OWiH80HnxHcuQ9L26IXDsLbbbQMViF6K+uQSxcxk4RwIDZFUqrCyQC1
BmDcmJ9jFbvigKHBOZXyDBzennhTPFGjhQQiPybcgQPe96HsODeH/FfYCM7Bfvih
oz4AZTnzdlRMU6ZQ7hOtMTkZEAusa6eEZ3SFtj2LYX94ogUvdc6V7s3oH+u/S9D+
nMTs5fjbNZrU/+tDdP2gw/sTwnN3FwbQJWyAljrQLxubCfMR+JX8oPFFLEzzI3HR
Kmy9DpTy2SG7DKt+90CN5cgSYUXprFGGHj+tjaDNoUOsR+WOtvufca+NJ41oWHGx
H6o9oHV/Xi9G1JftMO1AA5HSD4xf99oHJiacDNV+3s6vIn5ChkkEhgnyT96tgcUR
9UgF81rHpVt5srfW+eHtwhP8/Lq7mhUdxe4Gpv0OnqGlGsglwwcHvf3y82eXp4El
iZajmhejPnOqpkCXyu0mhORZ3TDrg0l6L8a5fKEcgomcD4Ep/7SLWdT8AS+mVCZe
j+3mwZSC3FnqY/76pJ7pcYuoEdV1aU7qOV6W2REIWEAs9ykOiYHzDlDCKrxpyW2W
YVAqXuLcB4yYVZzXhs1gIWNSGvRVODgkCxkVVxpXWPZfNXrmGJ7SRL/CXGloF7G6
Zh70ZZDR29aGxNwvJztjbZv9RUG4YdW4zH8kZdKrSwUkUUdhyMa3w0UJfTHHXDkB
4ddD9WRbuvrpDo20hmYHhl9pRIDLez7Yx9lRh2Sho34AHz2lg6tDUMPp9HemNtGy
BiJowsUoqyOrqnjyNuCwAbcwUlEZxiQ4w/0oEg+6EMuk9dCXIRqVhBklbbSQYZ2Z
SARowqGQpn7PhsUwvxIDQuuE02lgvetZVEviUge5pq8WZa4DySbgIUqyFhg+Abrm
dhEeARGyqkdiGtiLGpXR9oyuA3kOyTRxKtSpODGOuFjhewl3U9DF70y4mjQJV/YY
XCFSxljCFIgEIYY25etlNsi+smRvTFP/X3xnhqimROB7iDmVlxLGGil0FvZcSMSM
uQcWoJgBPB83cngwv/PbmKOtODTn0PhgHVKidJaxzGnEF6WdtYbrAAlWQdGi5ckl
5ugDyekmN5qX3smXRfglcYHWRvxsenxJ6RuHzrOF/31yjsn4NCKBfwF0OV3rdpDa
B5tm79LxBTRRPH2dOymzQjHdH5TJX/r8YgnhUM/v+qN1jK+g5wvr2l8Xk9afcbLf
Rfj6JFtVyeM8y8witwwQnwHZnxu+lQj23l5Xlruz+gBPpR7YvWXu2jOkCI6P40lL
QCHIfDi6ccYaIX8YXVgfpVGZ963X/a+kmxiIShtJaY7ptIKEC6frb16IoOhZhhx/
XnUmFsZIp0r7JYCy7Q44BmfBIre3jtgKcmO2mr0JzaG/Zq2qnx2Aef9vKRes/fi6
BWwhJhaDq1tdwWVl6Ic5GjRtGsjTu6kB+ovd35BIpAbeoNkOdxI/iSSKIyQpx1hi
0EWPOEosthjZGE19ZpBCBkEkBNuRvsSN07uy4xMoiRyitzsygQOA2iqqjNBVKXwI
WeDPxwjyOsLzs5XPVdfVfWoHJYIDOHforUldCYP9bpkCP/BVAPyylcBJFFNjKTsl
vxbNV46rsvv4SEVY9mYSniaM/pmzVh5hac1PEQXRzwxlYQS155lv1GJCch4CfhvL
7l25zR7kiQUBeAtomIDWPHoRFwUcmojZ422hgk7cOgMNeLq+sfPbFdvOwMiHN0Us
FWpM9mjkVeXe/PSi8u6W8XURH9J3ZfAjLPs9kkQny/8YuOe2TSlwWeZkGRg6DHV8
dpakV4l73xqgtfK3uGoiU/YOCny7gkPyCtznHR+uRlG5uQfVM6HMuipXg7LdrVC0
ebNzwR28sgGAnTwI+/n6GfzKYnLnLgJx9ojOvTdbNhHFFP1rDvfdVHXmgoAR9oUX
f4E8NaTTD9/AIW85E2cE5qrtN9jnoNIDlySsS/bN2MygNPOwFsTxnoaHOsZYko2t
5H3RfSh0FuyZ9ePg6qXEJsYoFeSCoGbRBpW09q/Y7ZQX4bpxNIVYCwkqW1yihBkB
5G/miXk05psYRVJA2+vcWFgD/XtaGH1DsIQ7Z7Gir7h2otFb15hJz2FbIv8NBlB7
mrtDSRVeviZdMWg4C3wWMloFQvKK8jWEhU/iU9HYzEyBFAkjoYkdZbslpvJT2x2i
cZymUCvNMKfeDjBT1Kne06pLjiSeEmWO7rw5KinLajswDlgoUOQqtKVxXw/+GPbQ
/xsotcq3L/ImKMAFpoyXg3Za3i2aSO0xejjOjHnEjm0Vj73SKqqb/5I70JOI2W8W
i0gTIv8Wp4tAPVkOm03VFw4wNlxNf6FSSDcewTZIHvYedh7M88BMeYtx11YA5gj/
Hpisi63n86pXebl3Ty1dYmUM+exX7nOF9FJ9XXhyjqW/1Rmb2kVw6541rSgDKV8y
a+mEdpVLZKKzTQGSqwlaivmIOAAvpXJ5eLroj/8XdwTSgzDyl2aw+G9EC7DjUfbz
1HUcfX532uWmpr+YUeQIneJFRDeMXu02CBRZTRkC501MnYt3qabP+i9j//Bw8G0+
AxKExUuVsfshgF7Phy0e9UFju/mDrS9SoHuIy6Yn74wOTRZrGJFWAj4zcygsaj4i
mAXkC05l4v2cDG5s6QNY64NEktOEwBBNu0HIGan11gzWzsuGLgDmpHXTpqeokvmH
AAnmP7YZbNzpQy/UT/A8KTQjJ6z5b7BbrEeCujYMgNvDvvLvK5uLOsrbjDXRiI8b
jZQlUBiwXGmRtO4agJPfZqUpgKqhVbX04Qtab3+2vPHT3rH5E3zGM5KuJpKXybQJ
ISclc1eVGsYD+Jzxx0jDIPzrdfjPVJYbU134PGfOHCzRN70PV8y/QTZZmK53pv+D
5UiTqHAW2TCizmZQme8h4zdaESSJ2a4Sm4BcuBgHaOo6IG7l6y1JXwhyCa1zyJsn
0fY55KQBd1q9EQ6HwIPnCZgq39FvubCgA31DNIXKEa/eck72b0x6QHDDOsayahTV
Ns+b5bwzjLOtqLJDmPYFqbnDrq9mCKY1vuOc12CjYcPYVz0sH/qtOHBJ7tpCFv0y
MvfLzgC9Q4yG2s2V2FlpzhD1ww/3n8891dk08ysFE29Q1/pA8gde45FsFFEGRe9/
ukhyvZpjCDA7vTMpm9wf6AhYrgx33azaqeuCOS3gCTZihJ25DxfM2ScLSg0a491b
CjBxgc7iGPbyBRCtxIKHBMn2Ki9nHW04WrB0xJEXqjz1bAMH7TGnApowU8e3OUoy
jji7cV38hjxQJAwy2RHm0PUEKYQVCmgQxakKnK95s0p9KM+sadSE9f9dxWqZ2R0A
etqZ2tdckWpwwCIIXhRv+ZY3EafJMwf7CzsCt7H3xXdRFMpj9gd8S5cfm84hZS+F
jaiNdmf6nflBlS4q9hkKzxy4U9/ifcwtbTTQZd7DOJ0kq/bkrydWhdF4yfJN1diK
hlK/WAZ2njDM4vbpqfnAM+QqfoC6PMsYlX7TSEnMoMiX16OG5HqQxtKMELMG5Y8y
oWCLZtPa8loRztglT8+/JnHlTWjcmVGKnL9fNrLyDdmGBQMRhIXxMxnl920vHV4c
1ddc0I+VssH27n/47xoXR8XGclJTLcl074BgYK/9FnRYQ6fZ6hhwcZa5HIy6ugIn
sAOdfol5wP7YJdlO5qapS/n+MGzrJd4Ylz00TJrURe+JLu+WCjGGv8a3a+uJ5dEv
Vy+LFmev99Q3iy0wGRwEDduSjc8/wRAxxoUIESvS4E2iSOdy1kbzvzWPJ3W7OdYS
0BnaWWImxh/Pl3aKWSSmoieMcs76CVoj6nBsaVZv0ZV12T0rQNFEYrwz8AKydAeZ
WS6Z4GcXAV94xpm/QjW76pREP8sTB2B9Ba2joTsS7H3g1Ao2TnT3oWfUOQ3/Tqy0
kVR5p34wdbQI/khqA9fQCXytVANC5V+RiSL1DI16a40e2CaJQaclG1Qm5Lq5VRfV
QB6WtuqpZVgoULSrzF9VQ7Zvlnyjz3sH9JwQj6FHu6mUdXAI/DdIidog+S0k4+JU
YfTxphQnnL095vgfXNmGD7cRv6RUk8Qznzt7zCfx/F4CGaK0GNwT3SmOahHb6fi1
5fIfV8vG41dxis7n22g+qwm83C+RqMWR8EoPsBuuVLITyv482bNIHbVXgRBN+T51
O2kZF0aZr3hvcSZR9rrdihSzDbCGP3njYoU9PP3Je0zDPtYJtDuK//vbQbn4BDbY
Swu2nSGfvr5sJ4IzAI4D+Dxa7wfs6N95c8hHa9E/Z/cmfENCzXCiaZ9Fr2H19wx9
3JB7Ku9K8m7VPaLTubEoZ9+QXuNZkuhDS+Hn3QsYJvfBYdzpvhpwqU8E75qmvJXD
l032QTQu5n0HNJoxIQHLMW4qv7Iat0yIf30CSY8YxBbtCHNmXTta4+YJOGgUbIPy
pO1K9QLn4H0jG4G5XK6Kp3/tq+M54VCgu/Wuy5BJFK0H8sqirre4wmvnNnLqcaPy
g/zYpldDDAhTDdtpK+T1jV0rtNQ0qWuMbkdAjgataWbO0cHGonnCPYcDyuKvdpu2
G631AeAVQBZr+CqegI01bXxK8G9yyEUlt3KBJL654aoLv2d5Ar4Nrw3amAaV8UEI
IJt78vkM6wjDFKMjbMWLJSkfmDlRnkXaSPm2MQLazOwPF5AnpAYtsPXgYGfxnfIR
mV077InT9Dwwn4Bg4uWTtifKl9XyK+JK707w1ESh+EBbeloL7/LXJ6QWul0jCkf/
jYef8J0bTO85FXhZuwKs462Nh18B2gTz0kYkvW/LByj6TGTDH6rjnMeTuzCJrp1i
0vIwmchd5DGQnxKHe+EeE8+hE+9uUHBKfmnwPz+hxds6C/D/X+GIAjDdrru7W3eG
tXN67WuExg2GTAGEut9n9KpfOssg7f4pLHiePGc3/MA3ujl8AZx9OMEh60daAq4t
p3eK+EIJ9r/IhgaT7xgh9xXW1aWheCHhu4DDfhxHQHF61nJ0BrTnJeODZXVaDn66
o23dgKFbXmcDHYgpaQ/L9lWpFUO6fxkJTLCabRgOKx97kk43ieszjIBgM0/aNDTg
NBM39TZNGZgCAmwolW+4VNv2EV+84lfVrjgqM0rRoNEXXLW0UHFCDYiVRcyJ/OCw
ma3l2v5lEp0qtHsR7P1oMbpikrQTp6Km0cEqASX9sgoxp35wbPbYWEj0dGpw1k+I
c9ZwmdeUQ81whi6HdZK0gXzD6ngpD/MPctfVUKxHUD1gGeHvDteS+cM32l4uHzur
1psbIAC1YUszQHZv1S5lmdfpe1dpfonYeLseSYUd7olTQS2KRrpTlJugwDbftyQv
2M3kSgEcJr/RWNC8ATdulGTAiAfwGe+14iJADZl+14uL4aS3/+RbVe4boBEjSwj1
HjG5KhL2yCppJnbR1p1HGZIQCmfDEinjyGnNGfRA9q/1xdtFjQFylK2f1N8YVV++
gKU53djNMA4ircRshdJk1dSZ2SmfWcIO94WQfK3oI5s1NvsP+KPuR+qtfTzAXoSs
Ek7OIzCQE6jWYKRQ7BLp83tVuihC2EOpFulhCkGPINV2vk6oxb2tZbdsGyynxeKW
X539rX5pI+VA+03iCOMO9Qm4f+vtSInRLt57kGDJyvTmHhu1PUWGzSmeltmNC3lK
yhcRiEBsyAxQh+jQ9VodPattY8wnv0YiXfKt0uyGtaZlvSuMTXe2i9b17CC48S0p
AnwWci6EQFgUdusCXzgKXZeMknhGgYecFvFk+hF+weB3JFegOGegLFA5Q4pQQKdh
7TQw9+9+09hR3bcuFC++KI9H2/mtbHZ9NoTDiYt6+694qbGlyPoPXiz2H1SLvC5f
+22Y+NYEgNtmoxZB8PuOYqkFaUnIunjeSoCPtKN5cbRrK7P4ztliAwmNsCBuhmJw
JAtuGt4E36cXcP9wnhqzOC1b5kW1XTC5qOosa2yrf6FpC4gceTQkDyqvC8hqVfsX
GkDZilPTBH+DP9fAPw7G4+DrKUM3PXYgd4kAHqqkV3DclQI9R0RnxEbnxCka41N1
otFHz6x+zHCY8cglGb6+f7NKtf4D+bBuKpHvLKy9v+LKpibyEUS8P12OALjybppP
yKul3TIMhmOJ1CljCzNzbd3NB91rHsK4VvORC+RTRsVdw4QLSyyma1ZKD6NNc4ve
g1I5EJcKMur24CowcSMWztEF5YmPl5Oa5zEzNmEA4bFde1rj2Asc/m0i9+mJhexR
/ieUkhmW0IjHlB4DePl6PWgM1MAIujf4iCmFDUpgcf7WdfaLz58lamAdMjnnGtra
fZuzhDYDl0NZ4a7s4zt49/KybH6sbBsH4okie51WFwZJZ4fDCxREr3oY9u5uQa/4
cLzDlBNWyBp9XdeyvjZ/YNS4mwz+AHfc2zRJVzose2MsXTOgBAtb9D10/mEzwBe6
Qf+A20IPtc6cOMrFxjaqv8S07czEXniGXxtnpkpCI6iyNA7lXcbAAbG5+6XJMEDP
7i8q+6Tl+Et29LoiLRlwanuE94jInKffsDJtzoWSSwWecOnn4Fign7CBC9Tlu0jc
DsWpDRqbBeCdvKu8iuVs6Zlm5bXRIwAN9OaIf/btorX4e3+F0y77jaz6xwrNi5mH
v1kgLCG49ZWEUxwd2aVtM4AggSGwU+eST72cMNOba086TPhq+vFFSqjnhNfzFXnV
HgDQAqM8ICcrsFmuttXGlE5uk6fwNRTi6VLvv5+EVEnrKEeP6LEUXFx2KVIcKZXb
KX1uzRq4/nQHq9jQ23u/T0Pj2vFtuZSmN19CaMqP9ielWSyyaNA2IQKc+mS+PYxB
5So9e48bryHGp996dRYiHmMemroxEroKHVlvWHlteh4anmnEeSDYX9kdlwbDU+1y
dmDLRPiqRS/aRiLeHT4Dc24l1wOoqdcW6SW7VuhXiqDO6fHFGUTefbwycK34qwGc
gH+LYbWDAWYfLHmmGUzeFHpGHS95NljYRpTfTY/JlEPCnAJMrEr5OZd8YD0EJgEc
/+1xYSq8q54pjnUnoBx3tlKONeA6m8dOyaHCQMAytvpCNDwBSxhdR/0tf4OEp7Ej
0o08ONIEq/gPXo66lFnvpazoPFefl6cSaCf/YcBj6LlJS7AjBW9/aMqEbxqjzQC/
jMLkPGIwg+EZlk41pozCN1uow4moJmjG1KkogYSVv3qayeNiRXIj0I6DX0PgHY/U
bIL/6qHJ7ePQSRaqK7eifjbm5tSkC6BAq676z3vV0XFiXp36u9HSlHkc9AFbp6Xv
YRNRYlpfvW9ZrFwyEFItsEZYGui1Wk04hBzKwXIKRBCEJHd08EmNhAF2Iya8/uj5
az1zIJYv7S3g+oEefvriD4lckO9puOBhtPOYoJxu+fA9/LgE241jTj65tZmWmUv+
wj5Dft8H/mW75umVHzvsMkuK4hoyxjH0uZ+QTT8gbHzOkTrB54ZJUtwZ1QtOtNk7
sV4WlzoL0gV3RzZi9AXj/eYw4YswYiLUYL3xpGvFk9jt7l9yinuklPx+cGu/lTeo
wU9wAcgHXvIjghsFQR8ZqOpsAaDpB+qjV4Jiq674S5Qb1inwmzwx6+eoZ8gzvuZ2
4H9L7rFuQVHSjsCU6Belf7nyFH9nQPIxEOUuG2D1v4Yei3pmaoq5SSJon4wZMuW8
gwXe95KAZtHYPtLn2KzcxvpcdZ3e+H1mJYBe64V1M38jGKGubNWG0WjaLtP+Fkfg
owWHm0T4a24899iGW7a4egySr/3qi8LYS9eP9ijZMBgKieZ3e/l4kzvynrPVArsx
bghHyipGph+0NhogxN8QKIh+ybLDcjI6adMd/7DHWohGspYfiY9bZv2iIbvsc3aG
pTcBqejTo7na8LN7BfhFrqA4PAV7Wh89J1NLuWBvfzecn6uc8koH184oVMLHZRJq
vL8M/Od4WafYy0Xs9VEtDNm/YFSey7sPpWE0I0GMpwo4BM+D8FFs6w/HyePtR6k5
+VZQV4+DNaRCNqx2NdKyGCM3aVZSm1EuZk5mg2ZQ1VgaZZR0pBZhUcddO/ZzfoOr
C+XQONZNPvcoyo2PvHeIZLI6AjGYgXaj9ombrVeUIwi8KVvOyJDeo3n40DGW8LXt
Xaxwj3608pEpQkNC8vZho2/X8BQGW9QzucHw6D8dT8ugA9DELLL+o1ejTXRe7mw3
yZvm6vwBWCaJCWbyB8gm2FX6PeN2ELDSWbz4D/ujPwY6XBdYxl0sSzijVtBGScys
UqgM3eD0wRF1Ox74K5hGiV8JikpXIUBsPGcGpfYGr3CB4J2ll2CP8Nl0famjZHTh
3o5R6g42R15EPCVbsB9Gb4HzE4VWsg/Kl55HYdOJPzCJavQzJI9Vj6sTpf3aoZmu
+tp+57CGeLVutiQ5C3wGt/TCdH5VXRGLYzYaHnYSR3NJ1EMrHATaFm/7yOt91kUJ
mPQnw5/bbL2ALgf8lQLSSugHfPzFr5bD2pZOdhq7uM3AJQcLcE854b8vpLhkJGTb
Ynuou9ti+qWo30yV3lCJyKm2lIRsdJBl0azloJmfLnWUWE3CtbpcIuRmwfy1aHjb
CIZsqivP634e2lCoDdQ3I6RsoHfXRvSKMXbsV9efH6CnhdUU79TDTrhUmuI0DfUe
lbMuVXa8s7JijDujE++iAFpw25g1JiN2oNV9N/nf+HpXtf5YpcsiuBegxOzmkU9M
MnfQ409GJrKYv6WbmVKtffXhxG/FgBJW7WvvFtFkHD+Utm4f5P4ajloIIhil8Y1L
uUllgMcmo/htyrD6fj1lq53wNdLn97y8mcLXZDJUV96fDpDok2cqUCfi3s9YpnFs
k75DHAg5OuQvC8SEVdYzoYZtInt9h2ZhfVX1XrGgHpWicnBWUaYl8vMEVH/YAzq+
raIRpronG6JvvMblAV2RCzp8iE13EprCBEJFiCXuP2PYxwCPSFv1ta3Ib4kACe/z
fttuupv3TImbJTBfiPl/K55eYy3rF5V0JMcoItUvDOaIoLWbMyizgILLZ1DxDvvr
UZRehdHwrMXVO/MwOKb0oP5HhZ1mOJDliRECRbVD58h+RPoFzqtmeqJeaIOs1hQW
uFMhx7QLiWJ2QkBL+oPjQ5CY7hfMzU2UOeSONNmEFKwsSCGfl3KcPMIa8qfbPN8f
RSjUcoY64JdDPkR/kXtZr/8l/VP4Vd9rfAgwOhsTMxoJBGBfJzQN1rdl3A7LA4F2
QfoWXB80aSBy9Rv40W5vd4W1601HM4f9e1sUiclwVp4Qfzt2t8JNkWieQ8r3Vhsi
vLoyN69gEmdhCywGPoqgTOIoHFPtpFgx7zEjkGrW8Mbu5kZX9zclyy0Fj9ptYfmO
f5vjfHxDOx7F/d8xVC6VGROltMBqkv4MrzrxoYnw8wRKi4ggw0aWtDbybdWKQhYw
15ikufvQ3Tyw2yH1VcLTOoOvgpmzhS/yUaV2zF2mNGwaAajI9ru3OexXyjoyzMJa
cVTfh/gk6ESCxrp3YhHf/a0CBRbDiUQN8LkrtdA+LR327f5Tu6Y0qxerZw4VPRVo
JVRSvS4voCs3nSeP8M7I8qFarpgZKDpL9w3hjSJlIrdzRR3XOyJvoUQD6VUWNEsS
/cRNV+gGhq3x0+UpHo5agVh5/0EGYdM12zM9E9OUy/ZN/JT3IB6Yp3Tbcdo39HHj
ISMnzfMo2Vh5SI3TCl8an0Uq3JUJkndvdFOIgET3eDfD/Nbk6RsMwugNmaMOc3Ca
1R0rKXUuiacWeSka1H/pM0OgLTr86slfcWLLZ6s5eu5pEj85AKcRLMKaTgNWF/Dt
y5jfH5OlBmorLwtI05tNZBIWVYt0Jl3k2NYRlv2nM3cOirPfsl+4tvdOr0PJxlLL
ptPum0s32+3kceVv/RDdWtYBheeopbvZrrhTSpiUENZ4ONf0/f5ui79Q36Jnerkp
eXlt63L29xsZoUeHjRx1HFgV2BhW1/O2ioAJxkgtWSAYc/0Vehg2cGb1AWG4q6D+
eDNH4FXbH9lHpE+XLiEGES878p4/B4AlhgC4il3jqG2amMR2iWdPm/k8TnncUa2T
7GnHawNY4rTk13QSmnUZyyaIjLEke+OUgp0Ay8mULYQ5s6hCaMtb8N/Hz+Lzu1zh
7e5CIIqDKgFRVkO+g5aRuGm6vYKawNZcjoBiq1ce9AEHWqPkMEHqlgD9aSnUANea
5ftXmjbSIC/wteAeuMCJitZn6g4XEGC3IqD8+mtKeBVrY2I3vJ4+8eLlJoHzATCB
0QiRgX2fZ44DEujXUdoFPtWzqzA4bEx9Ki3eSqExtGx02zBreo8pCCFuVTPzywyT
OPfUnjjUTKViR+wpqb12SAFWRb5n0mvcaTD9WMD6RWXn3RnKidX4oCyLk/N1bhcd
42UrxLZvOqpjBEblQrv246zXGZryBzvCOwCmDxJyemMA6YacJwTeE7EkGamtIb4k
/meH9htVYZAYk4jTeP2UB/0gaGYNYtun5w53iGJze7jzknEiQO4U3BjQJcNjb1s0
P8qqor+r4Cdb4u0Bhli7kqWmGvEV/r2hznbKOvLLJ3zFPUvbnP0zNGNidGIS9BJy
xgcprV1yBWBnXde6519zw5j/n/+z0dRszqQ72OpAn5pavfZNFXTL48pIqgmKDMQA
FNy0H6mb3GVJINOwkklb3ykWBDIyMMMVTlPswzSXajQ7xPp8A5pan2JXtfAHHPcq
ltZ9KLZfRObdUoDa7SwP0vDY7JLOY4zlfZdbk9yc7f202sj+5O+5IECIux2bgfet
W6pQX+8hF9oDgG2mjVHsRoHEImid+2VFNHz9lr+ihNxh4cH7jPaPMQ2Vk+k8cBX8
qv3S+GVvQBoUgikSt3hm8gUu+4V6iPNVXPjUwVMXHCz5TMHi5gd28LTSM0haGFVv
s8w4BM6Gi/dJ6OgH/F5EYz1hGFLvd6FX6IL4rmL85/M793OznI/UlqnkDMLy5xbg
HDmCQatxQYzyoWq961msVBF9s+BWeJZXXSpa0HVrtq+pB+5Us69bP+6y9CW3lDx/
h2wcUyHBBhasG7g4hAfqRECQsjKOA8YIuGADXnLKakRwDse+3OWLz7gqR0MHowew
P7paofNURJ0tVWXOkYXXQyfDrgxf65Olpw9iK6Gkf069xzYJIUXPL9rI0rgotgRS
EWR7pSFDhY4x8bIWkFzL0XdeAPtfM8sMkx0lk+mU+bZ6lAm/zMGzaYRtoG9WkVXj
pkgLkxT6Ix8cl+bRXqqne4SG8IGmmKUdAOIvuxtVTerGgj7wlW6acTg5r+/DUMbf
kXVGwyHW/zfNMTCXt8xljGRuAFw4M7/D2MwL0k/JBP3YIzbLstRBA1gmppIfUHRq
aQ2Jiek3p7RnaO/UMRNPPicADUMNDp2r128UKIGOvrG+sd3PygIgKgrxCGoM+mar
7MSGsGPTj+wUWPs8iW1kQ93mjmAeHBTfg1Vf0vT4ybvBwNClHA1gFPiAN8i/d38T
dVMsCywdrKvAfpMJpNXp4xkGlTFf75LlIWjvJhACmxHx3v6xxUpC8mjmU75Pk098
ohKKnO8Hx31GNCInzXl9lTSPXknHfs0u4fBaWzWP/g6BMZeFoG8gfNJnyD/FBKoF
CIJK46L8nMwYxsuUfSUCcxIgiW9rwSXTsgDlqIu4nYIgrszBZCn+sTt0AsHkt0qB
kqquM+NwgCJtNLfu/xQddhOdJPNqpIUYvW/yr8nwoE9462JN5Bc8k+zynb0i6XLV
tx6woDVrGIsi1oX+qkWhG4C0lGGaDCIVMJxYyr2qTUn3RRKK9OZXVW5ZehmD4BWc
I4NlS/QHKeNpiRfys6jTZP7HCBYIeHNQlETPKCM+w4Nry7dV8kbhy6onp/I6MNzL
zQcIsdd9o69Xy3U/dpuoF1DNeFWdk2m7YjV8q8PJLVPRLq2QAGFwtOT7Zp7/JyoJ
iLXJtGE/fXDmNKVVpnRBwOHYbZygeItqq+r/VDlZzVWgIp3MTVlcTVHonYlIpOZS
iDYuysJrY43W+dq7dRbh6SGiC0RHGoNrxtTCFydfHQqMCUXsf8sZro3li14MnrrI
bcpE+BdMxuUA4aI/8uBSs7nEQMaNjEYHRPemo+GfaZODoraIZnKStJ8QKDkzoN1j
NrFM9nsX15Vu2zWu8UcY5ntMXmB6HdSHCcpGiYbjo6LPQb/5Bl0hpHRhagdimEcs
fOoWEfar5M7I+RN23C+zJWONUKdPug/pV2/b3g+GoBeKQt3SBmgBItH+B7g53so9
j07+1Tcj57FA8AMMMzLpiajixQh1JxdmML32qNeNoq1tDOdGd+wzeUHB/SD30dUO
Fk8T+TkNqUGvC95Eblps6vk+wHYgN85w0fFXchtU/C5MPsuvpWHH8VrQd4DLFg+a
DonPy/swqfcRxxaiFYDyWmBjoZRsYL2f9zAg8sb53ajJnnI19V4TtBq6Vyy24uZK
flNzwgle5b52CeGoySx4tod7DUh9EvgOBdzGfGdrfeiF++PxMn7fpc2vBXGtQZwC
66ddCmjrgEkSKR7wcqOAR9gbhAcyEPP9Qu2hUJPyWWL5Qn4yP5MFCNg6h39k8B8d
TG3a+2/9f4U6KVVWmWjttgivsgf4Sxhsw5rqkWEwMdn/5kcsc35FS+G1cLRf4HQn
QhLcLlgRSr2EH6gvpHzDEzMkPu+Wxj2rvQ49qEuN6X6+Uo3kqecInT/EPadsUEkh
BbbiN2oezFDIaEbYqzLcvh1er8lWXSYmXdKhr7BSXDu2IK16sMQjfhZO66vkiuu8
WAO7E9wMkc5ymmzfe1x3AjQAlLjnxbiJ5eHszvk3DwbQkwHWAtSgUQv+A/QVCprM
Mpnef50GM8N79L2paQ9Fk83so/OF5Uryg93FNcclBYYY49XiNOc1CgIPhwdjpBl2
JI55eRCdFCyEuBVpMURO6l1X53/R6epeKGwAdaJEZefs/xzk9v5xTwL643Urzhhp
inft9B8NBb/JeeKEmALBwlRdIgHePuSaKc2g16cJ89xmX8fRL575x004+pFWr2UY
5jG+EI867adKqYBc1MkBndvWKPTDN3S2qBIahtYi57r+4cqT4oZzLxml6o4pSKYU
bHiTF1WPiBsPkArxWL3ErcxL7huQ1A2hldZBd+iM962XXCWfKeWpEhPngUrBg7bO
7Cy56sqpl1/XECe0H/TVJBoSHnibjmHFgsP5KRmqHBnbmuigrXdpbBFGx07+BoQE
Mf0GuTROHEtfbYXn4c1zi66X7v12/azBxMkRw4dTTOZMCYrj2hqAuuYXbxXqLwyV
xcVlFdmcqHO/K2ue+ZN1pvAuU7OE9V1qTsrckAn/a8EE8Jt4WI02roDveRP5Xo1y
Y9Q6a4kwn43SpHNa0gk2OVSFddQ44RdrljWzz5VlISjelQbNbC17tb4NFLA4zZ9Q
D0QnqsQKQOM3erTXsUvYferb7GQmuzJ/bb/FAZNJQ5xU6Hu2Rw2PInqLa2Dp3FwX
QlThThHdL1y1hHvR+Nwwf1EvX2RdCRflJS3xtNBT4C8uNyKIOM3ZS2TycbvazwM7
h8OtD8aY/eEHIf4U+0wu3BKZ645ls1QaaN91go6U6nuDSFMmoUKAVoERxFKbGN42
dJazeEcVab/odDXEFkcbDV9Eoe4EX3NZ1DsDuIuMm1iufJlB7AbRJUsel6dqF1ph
wgi3MbuwUIsvNlOuWcS0mS0VkMPFho5wbGP7eRKCPa4HjeKF+eXXvrH0gP56aWIv
muNB7p93ApuMJmJraT7656MAnQK1Y/9/y7zFpV4dTvkzkXWmT+PTj139I47+Mzb/
NpaO62Ix7NzPXEVM1UVjTs+NKRFlrdzev8JS4BtunuUsn/Lo1WHiiBcYDpLfyeXn
M6GvjW6YtoBUV7j/cJb5feS1OyM5XV36oOd+Rnl7N78GSrdQve4aGiuD2l3Of3dX
bZS0XxOaR2lPQMl4zwIksbKBAu59d3E08IwF50J6UPuDNADAtvPyKpPkCElTIJ09
Ltgt2acC63INlst3PjPkdrB3sK6thuwTPrLh/ktBWljzE7xpnOJ9XHBEcG16JfiN
fqS2Hp/03Vq+jVrViDaEn5qO8tL6V+ghidDBxXBFlaH59ffXAvKAiAiGnn37obrV
QLtbNLugSCxfVUvgiJl7LJfuoe4m3hi+W+l1PN/r/ozGLmv9XsYciG7idUdGb347
guiBA/Qc4RaQQTxGTfvoXAC91nzzdtl+u8mmYs2lzYRbQ2KecWu0xBNLwo3piTaE
iHC7676g1MV3Ik+9pw2vWD5ODKl8u/bpda273pB6gdWph/b7teHsbqBtnhAVXWvS
IpI+ZXvsvn5d4Eo1a4BkStAx/a5Ww1CaX4Wix0P0LxUY9o4v3Oh+mM2I9fPTQuTN
e6R0lTuVD+8Kxxmzln/g2D6m4+vKcFCSxIIm6/fZeF2GzvV81+oG98IwVwMH+Grs
+0jeBigQbZGE6vblxnVH755XHgnt9+lovdCmYNqjqMwOb/XlejQKXvkXZo2BOuIp
dnNdPkcF1rWeb4ir3RoD+VjgmVrplN40rWsDy9M2QZUWgUR7dMi/LT1AHXzJ8Jst
pP8Nj+jZ0RDYX/kaMnD98Rt8OE9iTTZfd6Fet5RvIJ4w/x0pDxuORZfec6WWElnl
PbVdrnlbynJoYpTcSRDLqBngfbulsBKyUpNP61/Q9DlBWPaILg7VkOzArWS6zvwb
41BP6Gb87O6IXMZey4iiiiSEzARoiMOM4p3xRrazF5jnCJY2kPsGIkdCCpVbLftC
SFLqsWVAtVBjYbwkODAiOiI2U7EgFH3HxOGdCKoc6jyFepuWsiNQE1G13IGakBY2
30+by8QnCVZoQnSv/koejCQFrFnngSEjQ671bw+sLbnPjWdMHei2/781Z4hpRoio
bx8lDzJHeZPU4H3dxzO/sEcxRU5vRWaXT7N15PtKoIUNpwK8S8H467It0XAGNNmb
TpW3E88D4q8blZSoW1DTGf3wjmD6NffOtpdZBwkkgrKenNkIGqYyt090LOPRN+TV
ClD47hDdilunTcSsQW6mK0ZfNQJ1sMvpVoJYUJvpDgGE5Jj+7PeGgUaT/f6HFKyx
/Ef37t2kMCtde20UybZce2CUFfSA3uW6G94W+/3EFqVt9UwdRfUNthCektv4L05F
FNVkM8R+R+GtnDi+ICCsGXtWN/LFZsQ2JGXSPfco7VvGFC2A2kD88a4Y0b2iuVFT
GHZHNVlY82R/ClheoT0I/LvyRcwgHAjIHGZa7yS2BUVGTnHpneZW36NN3kjx6pjh
ave5wEFUVy7LHrGZoXe50Sukl30qPnFUCOdZWzw+UaO7FmmKi/Bjl6pPAw58K+df
us4Q6L1HJlsO5JVgq9S+cHnyGlqwh47RDChKqfUlElgx0JaIghyH5Ls7sklxJUDs
ZPHhUHAtUe1GsGbNrJRT7jOGficXGfEy0bTW+Bx4vpIedrgMthSFrRymU9p7JzjK
HZbLIjUUz8MI5/xKw8CdcZqRrTvzivWlSxdrpELcjsrTXuMTlWVIiO1ki4C1r2C9
jzJoKAGsth3mV6bDTzcPKSh31qGtTuvFlQ7HEiN4YRCLRvq3CcRnn8Sugs6to4oB
3JPt1Bsxr/uoplZgANqGO6oSP56Zwbxdm6EEgWrbXP3jdJgj8c76ML38vqlchVQ8
/GH1D+mjYkG2hH/dH9J8LTSQoL4TsrZCHfb+1hhhokk9ZuhYHkgvIecLhkD52wxv
iJwSnkJ1Hb9uQh12lyERIPLdhXeNHRyloEGeIVGj6cE9Z9ISZPV7OGCJY8k5WvGb
86Cetqu1aRWmPDu6tPAs1gZx/Es7vzFs34j13CRf5s5pUPl/P3e86CJjWN+p/H+z
KtFugwqFpAep3N/g+zY06u0VCv88/u/YNW4oImyyBNZBmv0giEGYGjGQHXepOGBW
mOntWPMG/I9M9MoQ0Aq14T43we0WiBDiQ6kD8YdKka07acuc0JQUKfzdRQrqiOq/
Azg5gsiKUVqXvL25h0kbpCjmSFnu/XKmTJMLXK39h3AXMhvUIOaj7ZrgWhjxyq95
AIVK+PSCc4lkhqq3XPQfualNtizXbgDE6VpjekUZd2J5/MY01O382g7fIgXgzNAL
DMbIg8ADfg6TEaGVrQr9FST4uYu3Nf3ieAzRVfDb9xd4yCV4XAuXSHasCI5GJClf
H0w8hKnfo6+l/n7nyNnQqUPa4CrQ51vGf5QBW3R/Km55Co9P5oZsp6Nr/s67Rd8K
HADeWmDfCO6SXvcylLJNYyyCsMlEyrT1qBmODJCRQvuyWLAd3OTCNNKyopM8wJAw
yIKhxdUaclQECn0NllvzRk+kQLoItdUejtuoFTincEGttsZS4MlK6druSOyS9dQM
cOqeOXp9DzpHnDsn3gnkjEkurGZB7JAWXbKhzea+J6jRcsC3YBagz6hTPTGqqq+W
w72AoP5FgFKDO5yMS0DYNUPamdInNo4N5cDB7cfDRIlIP2Vtwh15oIG6lpAEPWRf
s7yAde+gK2P4JsQNmOvOxbvLILNBhThCInIApUICrfvCgWzcxkShv/5/yQds/IiA
aHTVm7MFm4aQ2wdz/L9v4TI4FnwdFDnoFSRlt+xLIf/iKWYXG4IAn3cf7CrsiZAd
sPA/ukD5PlyoOPGy5TjgoZ+1iVp7Eb/B2CEyhrYGObi96YzEzPC5wXDsdItFXUBM
aSdsItV9tMH5qpC5cYljmWM6DBkbeTIg8OCK3ET7dWaZO56hw60B2n81BcC7aa2z
PehJWH3B/OlQ8m46+2wctqpR+4wdpa72Lt9kMQxbNpvGPrq8PU04nzRzMmDOBteG
dRL3fC2yTO0KbFyjAoUr1fCeVEWfsNRV+9XJR3MwdQbviCju2RlXIGpK4czGO3Tu
h8Ts7C6i/Cv2NviU31lifWE3f5mSHLRamSSDuw4KCw8lQIfmWwXm10/XTKZoiQ7k
cPc3/Jji6EB2VnYvc+j2HkmvVcb3CVHcLTvKLF332xHCu41+/wT9VvK83ipVnNeF
e/1k9FXqF1Ao9zBa1CdIMklVqBMDz9Ekhh5bDEVn9hXIZfjOkvzsQIjS8LcdIcb8
iQt/hJLH42PzM1WMQxCNwuaPAgtYKG2k5z7bo7Te/iIBHYYBQY7WBXElhHx+dJHk
c4elpGss8zZKKyXDLWjJOal27x375VyfJJjMD8lMcaXcSUIHkY3hoe21Am7xTde4
qdYFN2HMUtcCr+gq9b+/Zeu858lsAgw5VYR99JFrE4PVgTsVuo+Tt7+l/Z1iZ5lq
xFZ9jZnS8G/u8C0+mDIeFtCx9hY80Lc7lTumUgjF8gef6frt3Av5z99VOZcNHQAd
gSGmj3U8ReuAz3ujLMpYcT+pMGR5fsbaYqD8GNkJ84LQIF/42jIlpFN17D/X0tPD
RLYFEpqV1i6X59mLd7tB1qtFqHn2osVvfq/F8SQ/WDcPD8tRIyLAM7AbX5yikZf7
SHtrM7RFlXShbJsBShfqa0g9AWbxaCLCRS4lOZa2JMNAcPrZHqzYy3T+ZnEwNaxN
GDWMO76Zd1egMmZuSTVC94nnusc4yxVZsM0izcvYfdQsjieBfgHF1FvML2OE5oY1
HkkxUaTqbLxx8vt8MRekKstaTFuQEDWoPM1MIJaYUKksHNSdr8nF5ygv7XY0hELI
BCQPT99Wm1qveNcgSOaGyTICYJDJPqZVfIeqaFt5Louzh/Y96HCTFAe146+cdtIE
7REPTUu4YGs/3pzfuMTIqV2lA8pPm8qlXT3fptCvVWGuCHSh5vMDW3WopjjUUwOr
N6341d8+ZdX/jw1ca0fjJnULjvDqv61vXEwJR4Aw6PkMZD5FewIiwCT4mDEMkSYb
orTZrfvJ23f22YjDRvuSjNSakBmW/PfTe+uvC6b6nw/JHewIEoRFj7cLKpHkfnYe
jDp0N/dEDM8N4y+XPwRL6Pdk0kvKISZSG3n07nGbbCDJFe1WZ5ez9FnGE89H12Km
z1+AUSwbkfiKTOfgltwLEVTiPq8y0rRTWBdYzJZpGIG+C76InsJ2kf7XFXjn8oFi
/LoivG5sRd8znDcM1Z7Pyor/oHM+hnGoPi7HI0E24zvnTQFB9tpxaPi4kvie2AjZ
Uy10qXn8Am5UGsxufQddab3QCnGwGphEScANmUdJvCP/QZ5oeuloN3f4aLVTlC3u
l9lK7I/uxu3679qDvVUdSf4mzyVF4nZdx4YirB8NYT4hXrfT9Ql/V9JnDp/fSiaa
UJSHe49rb7A1xYG3GnRR4lXO+mAu7oWK0S8oOgf3AhlOf2KmKopRnXB5NM80yw6r
jMGl5e76Mkkzp7gxR7JRyH9SJl7SmDi1iUdkyDpS63vOyNC34WC+9tKXdWsFIsGC
CvpqIiSkWFWSn9noRHZ4bPYwdCZQLyhw17f1dwpwONcxQr1SyMIw1+maOZGkEg2H
YRpKtrDlr+AGNSOKyewJFAfTjlw4cJraMGABi73jt7FneFzzfx/gIueUeSK36Ywq
nBjkl2XUfweswS2A4/a2jL0Mqucvw+EAqf+0y3mGme3IKOJeU/AL9TH4sCdZwPQC
bj6GUwVcDp3XKeoJf5zhqBlP2/e1GrSbv0z97xXQO0CWFE2VpFN3JDc+Ctv+HN5I
lwXNznlbSEPRFXJcz0d+6J6wphComGH3G5La8i0acZ6cX5+Wob9KpXvMcf4jx6Eb
E0O7yJh2G3tIe6b5/0v7IHzh+rrvrYnAl1h104T/J082SGi9JFh3dqX1HRTgezsB
GRO0BZowXeWA9kPA7/9CvD3abWkmf3KjURR4nM1QwNamLm9SNHjoX/QdfOGsRArD
AS+xILvmtMvKZ+NwNE30hxcMEj8995Ibo22xnUmij+ZgXRisiAEkHPDqjRpFgLbH
j52uwr20BHLH5OGXXDJMBxSdvuUcXWR5SB99XnCW+Y/v6mrMf4C2lzBV6wiv/4pu
nO+jo5n+oO4QCCEJoppkFJHX2B9Iu5jMCEhj1Yioev/WSbIGB4+cK05uxGQt+X4/
W2BeaKDhS9UiTKsi0zrzQb7TjYLvJd9fGV3HDF5jrJR7yV23FbHEXkB4eNuE8uJZ
7aasMvSATUx6fwihimvdOJVes1By52wbcPp87jfraBP5SXEcGCm1IlFKpb7hg6MI
EpXT20rXwo7yL/KF4Y9NKAqKMmvTE9+/CREdoFqneMrYXSmfB48r8s4dRdHGQn7A
9y4T6xPR6zNsoXTO3Q6AnKWPZm5N7+TFMbocJ6r6Sffi6mQCaDRj4mDoLeeUMZXg
Q9NSCWHbHZOzlXDs9yu44oO8rPz34cJj7cxS3YXyxu6TO6HjYATh9wB+QCoFpDiY
Vav69rZGK2qg3fonMw7kTqdPn0+8aiD4CK7MnrlJ53z0Tyc6XupY1jUS+BdtxEbU
/nxnZmitvTXdYq5LSx/8GEOsmfsWnIEMzivwrj253DyuzLl5nE+yUfyQqOh4M41M
1YLCQe+i1HSdBKwxQAr6rJPpr0FpEZJpYQAUMOsbqArY7WMj6xKIsxENGgc6Ih2U
xwcvBwmvsexlHnY5SWgh1gIEWUEn2T03RpgBx3g3y2vN7VPlNOVWIfNqmS//m4OJ
Xy2rTEQfsZLoC+wslReX8XQwiRKFqL3IqpuvbPhx7LTkvTcfzKQum5ScfZPMtYJk
6UgqFSL1SxlB8QcUu1R1fYnc1Vh6iJLVC5lWVjseaF3HizYHk6Yp0LlpqPpbV4N1
+H3YbvUMm9MXME/psWHOliYwSYaFfz+46DjwHvHFNU9qfBO3qKrieodG76WLco7b
a5ejU19zG4ei1XKEtdsvENXCaT0Kn+iN34qXAXKBzS4r+NPOnqOYYgPZupnBHdQI
CsremtC+G0Ho1ASpFbx9fkfI7iVAi5WNR8c6gGrSmEtagSRijNOTZSlmMQi6Eqto
CR4JbKi0kyaK8PcJjEhGVGMH8r2SsD4xCRZQ060pb/YxWYDkywuIqUR3Y4jhZ7e2
Gd/ZRlVJ5zoOJgvfYpqt/dgMzOJw78NV4zwbxcddHNxW/F1e/31s1fCSDj1VyADP
i4uub3vxdGBpJ4COgoMfCrcRmYEbasql+J8pplYpfYlzoP2SSVzzz4v3IlhoQTyy
gVmuAZ51mEHMxA9YgrOfyeXzEsiObFdE0EkibG6xVySuL33L3tuunnt52We6CgKE
GgDUN0wZNpftOtxwYQG9Bm5o6JeTj5FQz1DH2K1Hn4EC3rPQtt9bhACdBdlFkZjJ
f1X4sSp7adlJnpP58E6siITBK0Ypq/bxQ7/6QSzLzSOcfvpzpntRbtUZVrjW46DQ
hHL2TctSdRpzPVy8/tAskRB/lZ5z5bbcqpaUhCs3arvN0vymWEulYlNgFQtV6qZH
rPwdHIXcRy8aLtqRWkOf0sVF25TK0AeNay6V7EiBX/NyPw8IBocCpIMP0zCul9qh
vyTYg92cF7Oxs7aU7mzmOp0jIeoEPiu6ouTbYnmIYXSKCCAKGWn51K9UrRuxI0Gd
oY1wziEefn3/e5eOGSSMK23eNsOPb6iFYI0rRDtEbHYrJ4TSmWWiomm7bSxRCeDp
dk1YTFwZVd9Wug4bYzeuedYcxU9mKAq24ne8tdyAVAnUPaECDcFiM9+QubTInLi0
8mKn0EdCLDpV/kHgwcQ04k4ogJp23B20sFQUScODyctASk918VyyosdLxpz09DIp
H0kEniPGOVlKbi0f/E2Eupr7P7046v5PFHMeJKUGfzRiHRdZzDYYrmE50v4hJmAb
/qpsDmJ087FWyFYEBPaQs8z3C+Dj6LyTocpotILh1+70vkMLS+IqhKQ9TRXrC8ZG
p0KCbcEbomPmjfhR4qe395GJsOG31GhXJ09cvHeLpqQbHTauYOqdeQ1dHe6MdK4I
elCJDhV67Z7O0Le0ryaVAgLfOeIzwzKEFyqL+70ODHWeu6TIbLFvoGT84EmNP7ch
4enpkAO9I+ukBybRXZ7BUwpJYJ9yi+UzKS3CGrScf+m7jo3rmhELv1ukf2ud3DFa
rYdGsv8NTDQNN4pXn+MrkPzJQDTelS5I1atUeNeKRgYwMLyQbLea5jo+f8lra/Zv
LRTy8g+u4o1eADpZBQv5MfNg9FRq2c/h+wixE2INQhIgxIRx5btfF6AAuDcyhJWR
hUFSxWCHcAT4LDzFkIP7cZEV+Rvzk5EZpiRbqkCYcsKtYv8y90+wEf0AXW3oPaz9
vl/qv55/Q6BSV5zcqSG2MTBBm1h2PIBYDYizkpeApdL9Rc//Wdx6tBUYuhsiyFam
vHcQDE5Ch2BSJwSi6MZdsD2uLW2vMVB4AylW25XLrZk/Kq+hkWmT9Huu2wn5xKMb
zPy5Mv5Ui3uT1UKXmt6S1IBhT37YAq3N/AoutH1ePiyFoU/I9manGvQz3ShoJ2ZK
BUWlxaM+WD1tBmhyK4mSQg0Vocn13kZpLuuKFDA7SF/9AG+ZH9SofjlX7PoDRTVP
/4SAW48Gz9IGX2MXzkksu0Tq5tTAGreIs8BxndmKSwX6T+xrCRexm652uOrz/oBB
NQnXrElpNrKpyXRc6/wzPMyH6WOzDl/w2fbQLWTRZPnTH94kbXK85sLsyFl98f7c
Sxi91PneG3To2sQrK1H4zcDwzXrwVnQ1YW5JVuqb2psbDd5rh1Md7UHDWHxgW+KK
jEw+2L/CtwDlacOyUBARHpqPawJVJuv1Gy7SrC4itKIjRxfKxR1r5BFNSfAITB44
mwOopUv7Bfv589aD038neJKq4rRRYXS0AFi68HIT16h0YIZV5HFYDZRDugZvgajs
ksdahvqV6xrW+LD+c2mU7elbWBmc3AuYaICjCGPsY9COY+ylOY9HVE1W/Y+lZHpn
o73KN2dSUpQbxQbddG8NAif+pGFidKBvtUkt8f61CWLYiERzUfgQZyS/hFp+HcXT
uAFB4d9eYYvwILKSy2r0RqkZ2dUexeBtBasJCsUHP4xxOvFk1/ySVIt2Qf7os5JH
Cazknk00EFCK2HEk+4nOdh65vq6/sYTtWD/3ypPHKF/088KuoXgR+pHg9ZWQHzAW
sIr0yKZKURxea90+uhTdbG27DBTNl7EI53Pt4N1KoQdg8kBo1gMEArx2HyUtEmpj
SDBYKQ59Nzhb32ve58ezBRk+cI4g40o67Yyg49QhLRhjWPemWafgKGzJgqaoMIj0
FbiOInso5/pbvuwDX1F8P3qQyZ7eLmmDoaI+cSq+nNoOJtRo39T0Y+jkmRb5K+J1
+HHoSbpJpOsxMNGgJ9sxCJF50Ix9uA59aeGjAke7pA0XNqMqwT8ftY0I8S/AT01i
lOp40Svp/FOSK+WydSE1k7f0Fd678oIT5y7qreZKiJdvE7ElNdNKLDr4XfPrtHoP
nA8U6sEYxBTEsuaL+AIDYglCW0yHHzbDLOzGOJL/WoRrbT0x2Uq7OgBz8S3WkRZa
E8CK8p7RTzWfT8oaO5zh7Qx/CHGtU83eaDiLbhlnBAs+Tn+T+Oa7/c1E2DObNeCu
Z8DmDxKEQOhD5hE0HvPIxvUCtqHqpx+kPdK2zH+swnR2hbtj+scwqwTOjxCKjGJx
KuDzhW7ycBRb64NF16uyke0p8T1tQIqWmAE7Ogt/76LFAPbQNvPqnNLgjzJVnKeo
eIc4lR91el4+nXRaST8/kCxvfBk1ZgVbXbyk9W24MH/zaotVhQIxKfF8C1RsHdlk
4c0DEofQhZfQLYgX+EJts+BKFOVLGyVBUbNkHvUiRYjYU5oEuvTZ96yDW+hcUTKy
fqfQ1/ronvUwwanN9fFNKRsUP/y+eySOfMPAe7/sTTWO53gU/mX8Yy9BllBOomf2
tMhDCYVa47NF0PjJOyp4Cm+etCW9YGKkHO6bp2Jgw5ZJf5GpH1kMvhrs6NZbtexp
aeeITiO0bMHaUasXTtQo2nFaACHSbJCXdguD+QoTEwCxEpOtfxCBRbeeBRkbq/Uu
HKYBdqzvHD86cBzJj+KZw9CiEa4k6JeFCpHJ5S5hIyUaz335g8KWoLxzN53u6K0V
H4I2eNC1HC2KrbgC83mY2A==
`pragma protect end_protected


