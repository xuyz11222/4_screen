// Verilog netlist created by Tang Dynasty v5.6.71036
// Fri Sep 27 10:21:13 2024

`timescale 1ns / 1ps
module divider
  (
  clk,
  denominator,
  numerator,
  rst,
  start,
  done,
  quotient,
  remainder
  );

  input clk;
  input [20:0] denominator;
  input [20:0] numerator;
  input rst;
  input start;
  output done;
  output [20:0] quotient;
  output [20:0] remainder;

  parameter S_DEN = "UNSIGNED";
  parameter S_NUM = "SIGNED";
  parameter W_DEN = 21;
  parameter W_NUM = 21;
  // localparam W_CNT = 5;
  wire [4:0] al_1deac949;
  wire [4:0] al_d0dc52fd;
  wire [40:0] al_11033702;
  wire [40:0] al_1c1b24e7;
  wire [20:0] al_1315ed94;
  wire [20:0] al_9bfb1470;
  wire [40:0] al_248537e7;
  wire [31:0] al_563a08a7;
  wire [31:0] al_dd9da09a;
  wire [31:0] al_80e06344;
  wire [20:0] al_327525b3;
  wire [31:0] al_50fbc01b;
  wire [31:0] al_6e5e4cef;
  wire al_18e25363;
  wire al_496fff9b;
  wire al_244bf368;
  wire al_55b210dc;
  wire al_f39a7e9;
  wire al_9762a925;
  wire al_ef2ad0c3;
  wire al_e7f7dbb1;
  wire al_b1f223c3;
  wire al_e7086bfe;
  wire al_5e7e4908;
  wire al_d16993ed;
  wire al_ae0a6293;
  wire al_d07a623a;
  wire al_126bbf82;
  wire al_1aac3445;
  wire al_f5516224;
  wire al_91108e0e;
  wire al_a4e1781b;
  wire al_dc44be48;
  wire al_d8dd00e3;
  wire al_a0bad8f5;
  wire al_c93e73fa;
  wire al_6ea85cef;
  wire al_52616de9;
  wire al_114eba31;
  wire al_c61b4192;
  wire al_7c174651;
  wire al_e05a8afa;
  wire al_fc3ee0a5;
  wire al_429ad05d;
  wire al_974cade6;
  wire al_a7f61ab5;
  wire al_59ce2e47;
  wire al_f91768e5;
  wire al_8aaa10e2;
  wire al_eacba872;
  wire al_443ad4c3;
  wire al_280e82d4;
  wire al_e395b4b2;
  wire al_fa28ed9e;
  wire al_2ae86398;
  wire al_12bfe065;
  wire al_13513659;
  wire al_dd49840a;
  wire al_76bda18f;
  wire al_8b6c63fd;
  wire al_b751334b;
  wire al_ad866857;
  wire al_99deb495;
  wire al_2af0adaa;
  wire al_acc29700;
  wire al_9aeb978d;
  wire al_9728d08a;
  wire al_8fd594bc;
  wire al_909f7a83;
  wire al_4c67b15e;
  wire al_6a58ddd1;
  wire al_68c6af9c;
  wire al_20d542fe;
  wire al_b8a75adb;
  wire al_d52efb18;
  wire al_9a55ec0;
  wire al_dc502686;
  wire al_6df3b432;
  wire al_ee07af72;
  wire al_70a23447;
  wire al_39daa3b4;
  wire al_ee504525;
  wire al_6f06fbb5;
  wire al_5a39f5fc;
  wire al_d9e84cd9;
  wire al_da87d709;
  wire al_7710708d;
  wire al_7b53b30e;
  wire al_2146282f;
  wire al_3671c669;
  wire al_171a84f3;
  wire al_dcc86852;
  wire al_99c022aa;
  wire al_b48babe5;
  wire al_2b1244ed;
  wire al_b54e7dc3;
  wire al_47b10981;
  wire al_b32069f9;
  wire al_60f185cd;
  wire al_eaa7ce0;
  wire al_f69c20e6;
  wire al_5812f805;
  wire al_a3d21b00;
  wire al_b2a0a3a;
  wire al_ad38578c;
  wire al_e110622d;
  wire al_a93ceae5;
  wire al_f2884563;
  wire al_f43e2390;
  wire al_9b8feb22;
  wire al_80ba6c2b;
  wire al_f752ffb3;
  wire al_30ecd40b;
  wire al_547478b7;
  wire al_a0f967e6;
  wire al_a629ebb4;
  wire al_3f9c0f6c;
  wire al_2105c1a;
  wire al_ec383fcc;
  wire al_a24ece81;
  wire al_ff12c8b;
  wire al_ad33515c;
  wire al_d4dcd819;
  wire al_d69530ee;
  wire al_6c403517;
  wire al_754ea4fe;
  wire al_37bc7186;
  wire al_2219a139;
  wire al_cb2a582d;
  wire al_65ae4a67;
  wire al_5d4ddebc;
  wire al_d5e7ffcc;
  wire al_a8ba9585;
  wire al_e7839166;
  wire al_73979547;
  wire al_e60b4bec;
  wire al_41c40f55;
  wire al_12148bf7;
  wire al_62db1d79;
  wire al_c5cd324b;
  wire al_be189310;
  wire al_a46328dc;
  wire al_60559583;
  wire al_c8377ec7;
  wire al_e18beeda;
  wire al_3827637d;
  wire al_91f93bf1;
  wire al_c0ec79fe;
  wire al_e662d6df;
  wire al_2666c71d;
  wire al_1f2fd634;
  wire al_f1a38dd5;
  wire al_4ad78cf7;

  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_ee4dca6a (
    .a(1'b0),
    .o({al_ad866857,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c820716d (
    .a(1'b0),
    .b(al_327525b3[0]),
    .c(al_ad866857),
    .o({al_99deb495,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_821d2ac7 (
    .a(1'b0),
    .b(al_327525b3[1]),
    .c(al_99deb495),
    .o({al_2af0adaa,al_80e06344[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1eb6e7f4 (
    .a(1'b0),
    .b(al_327525b3[2]),
    .c(al_2af0adaa),
    .o({al_acc29700,al_80e06344[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5070be8a (
    .a(1'b0),
    .b(al_327525b3[3]),
    .c(al_acc29700),
    .o({al_9aeb978d,al_80e06344[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_199b9a22 (
    .a(1'b0),
    .b(al_327525b3[4]),
    .c(al_9aeb978d),
    .o({al_9728d08a,al_80e06344[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_194c9640 (
    .a(1'b0),
    .b(al_327525b3[5]),
    .c(al_9728d08a),
    .o({al_8fd594bc,al_80e06344[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3fe0a249 (
    .a(1'b0),
    .b(al_327525b3[6]),
    .c(al_8fd594bc),
    .o({al_909f7a83,al_80e06344[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3d75bc27 (
    .a(1'b0),
    .b(al_327525b3[7]),
    .c(al_909f7a83),
    .o({al_4c67b15e,al_80e06344[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ad639e (
    .a(1'b0),
    .b(al_327525b3[8]),
    .c(al_4c67b15e),
    .o({al_6a58ddd1,al_80e06344[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aede42cd (
    .a(1'b0),
    .b(al_327525b3[9]),
    .c(al_6a58ddd1),
    .o({al_68c6af9c,al_80e06344[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1252e212 (
    .a(1'b0),
    .b(al_327525b3[10]),
    .c(al_68c6af9c),
    .o({al_20d542fe,al_80e06344[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_802d6d3e (
    .a(1'b0),
    .b(al_327525b3[11]),
    .c(al_20d542fe),
    .o({al_b8a75adb,al_80e06344[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1f07c543 (
    .a(1'b0),
    .b(al_327525b3[12]),
    .c(al_b8a75adb),
    .o({al_d52efb18,al_80e06344[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_50fd806a (
    .a(1'b0),
    .b(al_327525b3[13]),
    .c(al_d52efb18),
    .o({al_9a55ec0,al_80e06344[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5eea9400 (
    .a(1'b0),
    .b(al_327525b3[14]),
    .c(al_9a55ec0),
    .o({al_dc502686,al_80e06344[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1d94888c (
    .a(1'b0),
    .b(al_327525b3[15]),
    .c(al_dc502686),
    .o({al_6df3b432,al_80e06344[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_69249942 (
    .a(1'b0),
    .b(al_327525b3[16]),
    .c(al_6df3b432),
    .o({al_ee07af72,al_80e06344[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_182c8acf (
    .a(1'b0),
    .b(al_327525b3[17]),
    .c(al_ee07af72),
    .o({al_70a23447,al_80e06344[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f5bb9d7a (
    .a(1'b0),
    .b(al_327525b3[18]),
    .c(al_70a23447),
    .o({al_39daa3b4,al_80e06344[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b8aec0d5 (
    .a(1'b0),
    .b(al_327525b3[19]),
    .c(al_39daa3b4),
    .o({al_ee504525,al_80e06344[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4d29a2f9 (
    .a(1'b0),
    .b(al_327525b3[20]),
    .c(al_ee504525),
    .o({open_n4,al_80e06344[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_d7adc91c (
    .a(1'b0),
    .o({al_6f06fbb5,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7f5bc3db (
    .a(1'b0),
    .b(al_1315ed94[0]),
    .c(al_6f06fbb5),
    .o({al_5a39f5fc,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7c0aa686 (
    .a(1'b0),
    .b(al_1315ed94[1]),
    .c(al_5a39f5fc),
    .o({al_d9e84cd9,al_6e5e4cef[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ba4c16ec (
    .a(1'b0),
    .b(al_1315ed94[2]),
    .c(al_d9e84cd9),
    .o({al_da87d709,al_6e5e4cef[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7682569a (
    .a(1'b0),
    .b(al_1315ed94[3]),
    .c(al_da87d709),
    .o({al_7710708d,al_6e5e4cef[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3436ba98 (
    .a(1'b0),
    .b(al_1315ed94[4]),
    .c(al_7710708d),
    .o({al_7b53b30e,al_6e5e4cef[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_91001818 (
    .a(1'b0),
    .b(al_1315ed94[5]),
    .c(al_7b53b30e),
    .o({al_2146282f,al_6e5e4cef[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8988f540 (
    .a(1'b0),
    .b(al_1315ed94[6]),
    .c(al_2146282f),
    .o({al_3671c669,al_6e5e4cef[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_66648be7 (
    .a(1'b0),
    .b(al_1315ed94[7]),
    .c(al_3671c669),
    .o({al_171a84f3,al_6e5e4cef[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6caaa7d2 (
    .a(1'b0),
    .b(al_1315ed94[8]),
    .c(al_171a84f3),
    .o({al_dcc86852,al_6e5e4cef[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_22cd0657 (
    .a(1'b0),
    .b(al_1315ed94[9]),
    .c(al_dcc86852),
    .o({al_99c022aa,al_6e5e4cef[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_10c9d72a (
    .a(1'b0),
    .b(al_1315ed94[10]),
    .c(al_99c022aa),
    .o({al_b48babe5,al_6e5e4cef[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d3583073 (
    .a(1'b0),
    .b(al_1315ed94[11]),
    .c(al_b48babe5),
    .o({al_2b1244ed,al_6e5e4cef[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ffd0770c (
    .a(1'b0),
    .b(al_1315ed94[12]),
    .c(al_2b1244ed),
    .o({al_b54e7dc3,al_6e5e4cef[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c1421b1 (
    .a(1'b0),
    .b(al_1315ed94[13]),
    .c(al_b54e7dc3),
    .o({al_47b10981,al_6e5e4cef[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_42b4a134 (
    .a(1'b0),
    .b(al_1315ed94[14]),
    .c(al_47b10981),
    .o({al_b32069f9,al_6e5e4cef[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_693341e (
    .a(1'b0),
    .b(al_1315ed94[15]),
    .c(al_b32069f9),
    .o({al_60f185cd,al_6e5e4cef[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b25e204 (
    .a(1'b0),
    .b(al_1315ed94[16]),
    .c(al_60f185cd),
    .o({al_eaa7ce0,al_6e5e4cef[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2854f5f6 (
    .a(1'b0),
    .b(al_1315ed94[17]),
    .c(al_eaa7ce0),
    .o({al_f69c20e6,al_6e5e4cef[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4cda9604 (
    .a(1'b0),
    .b(al_1315ed94[18]),
    .c(al_f69c20e6),
    .o({al_5812f805,al_6e5e4cef[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bcaa6e3a (
    .a(1'b0),
    .b(al_1315ed94[19]),
    .c(al_5812f805),
    .o({al_a3d21b00,al_6e5e4cef[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4eb57d16 (
    .a(1'b0),
    .b(al_1315ed94[20]),
    .c(al_a3d21b00),
    .o({open_n9,al_6e5e4cef[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_1ad5c4da (
    .a(1'b0),
    .o({al_7c174651,open_n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e223572 (
    .a(1'b0),
    .b(numerator[0]),
    .c(al_7c174651),
    .o({al_e05a8afa,open_n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eb751045 (
    .a(1'b0),
    .b(numerator[1]),
    .c(al_e05a8afa),
    .o({al_fc3ee0a5,al_563a08a7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_570fbb37 (
    .a(1'b0),
    .b(numerator[2]),
    .c(al_fc3ee0a5),
    .o({al_429ad05d,al_563a08a7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_49f69bac (
    .a(1'b0),
    .b(numerator[3]),
    .c(al_429ad05d),
    .o({al_974cade6,al_563a08a7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_be12ed41 (
    .a(1'b0),
    .b(numerator[4]),
    .c(al_974cade6),
    .o({al_a7f61ab5,al_563a08a7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1ab41e54 (
    .a(1'b0),
    .b(numerator[5]),
    .c(al_a7f61ab5),
    .o({al_59ce2e47,al_563a08a7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_efabd020 (
    .a(1'b0),
    .b(numerator[6]),
    .c(al_59ce2e47),
    .o({al_f91768e5,al_563a08a7[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a789b25c (
    .a(1'b0),
    .b(numerator[7]),
    .c(al_f91768e5),
    .o({al_8aaa10e2,al_563a08a7[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3f49f5d6 (
    .a(1'b0),
    .b(numerator[8]),
    .c(al_8aaa10e2),
    .o({al_eacba872,al_563a08a7[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27e18662 (
    .a(1'b0),
    .b(numerator[9]),
    .c(al_eacba872),
    .o({al_443ad4c3,al_563a08a7[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b30a8b98 (
    .a(1'b0),
    .b(numerator[10]),
    .c(al_443ad4c3),
    .o({al_280e82d4,al_563a08a7[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4f17b61 (
    .a(1'b0),
    .b(numerator[11]),
    .c(al_280e82d4),
    .o({al_e395b4b2,al_563a08a7[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_91fb82ac (
    .a(1'b0),
    .b(numerator[12]),
    .c(al_e395b4b2),
    .o({al_fa28ed9e,al_563a08a7[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fb284d76 (
    .a(1'b0),
    .b(numerator[13]),
    .c(al_fa28ed9e),
    .o({al_2ae86398,al_563a08a7[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dcc99eed (
    .a(1'b0),
    .b(numerator[14]),
    .c(al_2ae86398),
    .o({al_12bfe065,al_563a08a7[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_62a6219c (
    .a(1'b0),
    .b(numerator[15]),
    .c(al_12bfe065),
    .o({al_13513659,al_563a08a7[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d24a4ba9 (
    .a(1'b0),
    .b(numerator[16]),
    .c(al_13513659),
    .o({al_dd49840a,al_563a08a7[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5751e2fa (
    .a(1'b0),
    .b(numerator[17]),
    .c(al_dd49840a),
    .o({al_76bda18f,al_563a08a7[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a7bae841 (
    .a(1'b0),
    .b(numerator[18]),
    .c(al_76bda18f),
    .o({al_8b6c63fd,al_563a08a7[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a41fb992 (
    .a(1'b0),
    .b(numerator[19]),
    .c(al_8b6c63fd),
    .o({al_b751334b,al_563a08a7[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7c9c9a92 (
    .a(1'b0),
    .b(numerator[20]),
    .c(al_b751334b),
    .o({open_n14,al_563a08a7[20]}));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(~B*~(~E*(~(C)*~(D)*~(F)+C*D*F))))"),
    .INIT(64'hbbbbabbbbbbbbbba))
    al_f17cd423 (
    .a(start),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .e(al_1deac949[3]),
    .f(al_1deac949[4]),
    .o(al_d0dc52fd[0]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*(D@C))"),
    .INIT(16'h0110))
    al_147e6a1b (
    .a(al_114eba31),
    .b(start),
    .c(al_1deac949[0]),
    .d(al_1deac949[1]),
    .o(al_d0dc52fd[1]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*~A)"),
    .INIT(32'h00400000))
    al_c8620855 (
    .a(al_1deac949[0]),
    .b(al_1deac949[1]),
    .c(al_1deac949[2]),
    .d(al_1deac949[3]),
    .e(al_1deac949[4]),
    .o(al_114eba31));
  AL_MAP_LUT5 #(
    .EQN("(~B*~A*(E@(D*C)))"),
    .INIT(32'h01111000))
    al_56322a5c (
    .a(al_114eba31),
    .b(start),
    .c(al_1deac949[0]),
    .d(al_1deac949[1]),
    .e(al_1deac949[2]),
    .o(al_d0dc52fd[2]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(E@(D*C*B)))"),
    .INIT(32'h15554000))
    al_6614de08 (
    .a(start),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .e(al_1deac949[3]),
    .o(al_d0dc52fd[3]));
  AL_MAP_LUT6 #(
    .EQN("(~A*(B*(D*C)*E*~(F)+~(B)*~((D*C))*~(E)*F+B*~((D*C))*~(E)*F+B*(D*C)*~(E)*F+~(B)*~((D*C))*E*F+B*~((D*C))*E*F+~(B)*(D*C)*E*F))"),
    .INIT(64'h1555455540000000))
    al_6dc5f615 (
    .a(start),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .e(al_1deac949[3]),
    .f(al_1deac949[4]),
    .o(al_d0dc52fd[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b1b9ffd0 (
    .a(denominator[0]),
    .b(start),
    .c(al_11033702[21]),
    .o(al_1c1b24e7[20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b2cd7517 (
    .a(denominator[1]),
    .b(start),
    .c(al_11033702[22]),
    .o(al_1c1b24e7[21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e0f50da5 (
    .a(denominator[2]),
    .b(start),
    .c(al_11033702[23]),
    .o(al_1c1b24e7[22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f95f5f0d (
    .a(denominator[3]),
    .b(start),
    .c(al_11033702[24]),
    .o(al_1c1b24e7[23]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_12928f03 (
    .a(denominator[4]),
    .b(start),
    .c(al_11033702[25]),
    .o(al_1c1b24e7[24]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_2d4b49b3 (
    .a(denominator[5]),
    .b(start),
    .c(al_11033702[26]),
    .o(al_1c1b24e7[25]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_cdf87825 (
    .a(denominator[6]),
    .b(start),
    .c(al_11033702[27]),
    .o(al_1c1b24e7[26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e6264f31 (
    .a(denominator[7]),
    .b(start),
    .c(al_11033702[28]),
    .o(al_1c1b24e7[27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_934b4c16 (
    .a(denominator[8]),
    .b(start),
    .c(al_11033702[29]),
    .o(al_1c1b24e7[28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_9fe68c39 (
    .a(denominator[9]),
    .b(start),
    .c(al_11033702[30]),
    .o(al_1c1b24e7[29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_41104578 (
    .a(denominator[10]),
    .b(start),
    .c(al_11033702[31]),
    .o(al_1c1b24e7[30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_12c43e12 (
    .a(denominator[11]),
    .b(start),
    .c(al_11033702[32]),
    .o(al_1c1b24e7[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_ded93226 (
    .a(denominator[12]),
    .b(start),
    .c(al_11033702[33]),
    .o(al_1c1b24e7[32]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_c35e0dcc (
    .a(denominator[13]),
    .b(start),
    .c(al_11033702[34]),
    .o(al_1c1b24e7[33]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_362a2d70 (
    .a(denominator[14]),
    .b(start),
    .c(al_11033702[35]),
    .o(al_1c1b24e7[34]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_619d59f3 (
    .a(denominator[15]),
    .b(start),
    .c(al_11033702[36]),
    .o(al_1c1b24e7[35]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8b9da26a (
    .a(denominator[16]),
    .b(start),
    .c(al_11033702[37]),
    .o(al_1c1b24e7[36]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_14645c1e (
    .a(denominator[17]),
    .b(start),
    .c(al_11033702[38]),
    .o(al_1c1b24e7[37]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_41e73ba7 (
    .a(denominator[18]),
    .b(start),
    .c(al_11033702[39]),
    .o(al_1c1b24e7[38]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1a059b5b (
    .a(denominator[19]),
    .b(start),
    .c(al_11033702[40]),
    .o(al_1c1b24e7[39]));
  AL_DFF_0 al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_114eba31),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_affc23c8 (
    .a(al_c61b4192),
    .b(numerator[0]),
    .c(start),
    .d(al_1315ed94[0]),
    .e(al_248537e7[0]),
    .o(al_9bfb1470[0]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_7e4247d5 (
    .a(numerator[20]),
    .b(numerator[10]),
    .c(al_563a08a7[10]),
    .o(al_a46328dc));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_543ba616 (
    .a(al_c61b4192),
    .b(al_a46328dc),
    .c(start),
    .d(al_1315ed94[10]),
    .e(al_248537e7[10]),
    .o(al_9bfb1470[10]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_8f76e334 (
    .a(numerator[20]),
    .b(numerator[11]),
    .c(al_563a08a7[11]),
    .o(al_be189310));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_aef23a0d (
    .a(al_c61b4192),
    .b(al_be189310),
    .c(start),
    .d(al_1315ed94[11]),
    .e(al_248537e7[11]),
    .o(al_9bfb1470[11]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_43c29c9e (
    .a(numerator[20]),
    .b(numerator[12]),
    .c(al_563a08a7[12]),
    .o(al_c5cd324b));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_18f76fe4 (
    .a(al_c61b4192),
    .b(al_c5cd324b),
    .c(start),
    .d(al_1315ed94[12]),
    .e(al_248537e7[12]),
    .o(al_9bfb1470[12]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_dcb75b0 (
    .a(numerator[20]),
    .b(numerator[13]),
    .c(al_563a08a7[13]),
    .o(al_62db1d79));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_42d84427 (
    .a(al_c61b4192),
    .b(al_62db1d79),
    .c(start),
    .d(al_1315ed94[13]),
    .e(al_248537e7[13]),
    .o(al_9bfb1470[13]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_e1773c9b (
    .a(numerator[20]),
    .b(numerator[14]),
    .c(al_563a08a7[14]),
    .o(al_12148bf7));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_21d7d0c9 (
    .a(al_c61b4192),
    .b(al_12148bf7),
    .c(start),
    .d(al_1315ed94[14]),
    .e(al_248537e7[14]),
    .o(al_9bfb1470[14]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_8e3693cb (
    .a(numerator[20]),
    .b(numerator[15]),
    .c(al_563a08a7[15]),
    .o(al_41c40f55));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_ddb1c774 (
    .a(al_c61b4192),
    .b(al_41c40f55),
    .c(start),
    .d(al_1315ed94[15]),
    .e(al_248537e7[15]),
    .o(al_9bfb1470[15]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_79948be9 (
    .a(numerator[20]),
    .b(numerator[16]),
    .c(al_563a08a7[16]),
    .o(al_e60b4bec));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_276c7449 (
    .a(al_c61b4192),
    .b(al_e60b4bec),
    .c(start),
    .d(al_1315ed94[16]),
    .e(al_248537e7[16]),
    .o(al_9bfb1470[16]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_cd0015f2 (
    .a(numerator[20]),
    .b(numerator[17]),
    .c(al_563a08a7[17]),
    .o(al_73979547));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_d6e68fef (
    .a(al_c61b4192),
    .b(al_73979547),
    .c(start),
    .d(al_1315ed94[17]),
    .e(al_248537e7[17]),
    .o(al_9bfb1470[17]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_5eba52cf (
    .a(numerator[20]),
    .b(numerator[18]),
    .c(al_563a08a7[18]),
    .o(al_e7839166));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_754b9a1c (
    .a(al_c61b4192),
    .b(al_e7839166),
    .c(start),
    .d(al_1315ed94[18]),
    .e(al_248537e7[18]),
    .o(al_9bfb1470[18]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_fd435063 (
    .a(al_11033702[23]),
    .b(al_11033702[24]),
    .c(al_11033702[25]),
    .d(al_11033702[26]),
    .o(al_b2a0a3a));
  AL_MAP_LUT6 #(
    .EQN("(~B*~A*~(~F*D)*~(~E*C))"),
    .INIT(64'h1111010100110001))
    al_39e6fc26 (
    .a(al_a93ceae5),
    .b(al_f2884563),
    .c(al_11033702[17]),
    .d(al_11033702[18]),
    .e(al_1315ed94[17]),
    .f(al_1315ed94[18]),
    .o(al_f43e2390));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_eb7a60e8 (
    .a(al_11033702[12]),
    .b(al_1315ed94[12]),
    .o(al_496fff9b));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d22d973b (
    .a(al_11033702[15]),
    .b(al_1315ed94[15]),
    .o(al_9b8feb22));
  AL_MAP_LUT6 #(
    .EQN("(~B*(~(A)*~(C)*~(D)*~(E)*~(F)+~(A)*C*~(D)*~(E)*~(F)+A*C*~(D)*~(E)*~(F)+~(A)*~(C)*D*~(E)*~(F)+A*~(C)*D*~(E)*~(F)+~(A)*C*D*~(E)*~(F)+A*C*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+~(A)*~(C)*D*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*D*E*~(F)+~(A)*~(C)*D*~(E)*F+~(A)*C*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*D*E*F))"),
    .INIT(64'h1000310033103331))
    al_a510a139 (
    .a(al_496fff9b),
    .b(al_9b8feb22),
    .c(al_11033702[13]),
    .d(al_11033702[14]),
    .e(al_1315ed94[13]),
    .f(al_1315ed94[14]),
    .o(al_80ba6c2b));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((D*~A))*~(E)*~(F)+B*~(C)*~((D*~A))*~(E)*~(F)+~(B)*C*~((D*~A))*~(E)*~(F)+B*C*~((D*~A))*~(E)*~(F)+B*~(C)*(D*~A)*~(E)*~(F)+~(B)*C*(D*~A)*~(E)*~(F)+B*C*(D*~A)*~(E)*~(F)+B*~(C)*~((D*~A))*E*~(F)+~(B)*C*~((D*~A))*E*~(F)+B*C*~((D*~A))*E*~(F)+~(B)*C*(D*~A)*E*~(F)+B*C*(D*~A)*E*~(F)+~(B)*C*~((D*~A))*~(E)*F+B*C*~((D*~A))*~(E)*F+B*C*(D*~A)*~(E)*F+B*C*~((D*~A))*E*F)"),
    .INIT(64'h80c0e0f0f8fcfeff))
    al_afa39603 (
    .a(al_11033702[16]),
    .b(al_11033702[17]),
    .c(al_11033702[18]),
    .d(al_1315ed94[16]),
    .e(al_1315ed94[17]),
    .f(al_1315ed94[18]),
    .o(al_f752ffb3));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_1794dfbe (
    .a(al_11033702[12]),
    .b(al_11033702[13]),
    .c(al_11033702[14]),
    .d(al_1315ed94[12]),
    .e(al_1315ed94[13]),
    .f(al_1315ed94[14]),
    .o(al_30ecd40b));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_4f98d945 (
    .a(al_11033702[17]),
    .b(al_11033702[18]),
    .c(al_1315ed94[17]),
    .d(al_1315ed94[18]),
    .o(al_547478b7));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_6443e46b (
    .a(al_547478b7),
    .b(al_11033702[15]),
    .c(al_11033702[16]),
    .d(al_1315ed94[15]),
    .e(al_1315ed94[16]),
    .o(al_a0f967e6));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(F@D)*~(E@C))"),
    .INIT(64'h8000080000800008))
    al_49ff4809 (
    .a(al_30ecd40b),
    .b(al_547478b7),
    .c(al_11033702[15]),
    .d(al_11033702[16]),
    .e(al_1315ed94[15]),
    .f(al_1315ed94[16]),
    .o(al_a629ebb4));
  AL_MAP_LUT5 #(
    .EQN("(B*~(E*~A*~(~D*C)))"),
    .INIT(32'h88c8cccc))
    al_22a37a68 (
    .a(al_a629ebb4),
    .b(al_e110622d),
    .c(al_f43e2390),
    .d(al_80ba6c2b),
    .e(al_f752ffb3),
    .o(al_3f9c0f6c));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_304d7ff (
    .a(al_11033702[19]),
    .b(al_11033702[20]),
    .c(al_1315ed94[19]),
    .d(al_1315ed94[20]),
    .o(al_ad38578c));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cc178bb3 (
    .a(al_11033702[10]),
    .b(al_1315ed94[10]),
    .o(al_2105c1a));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_773b0bf (
    .a(al_11033702[10]),
    .b(al_1315ed94[10]),
    .o(al_ec383fcc));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_11a677d (
    .a(al_11033702[6]),
    .b(al_11033702[7]),
    .c(al_11033702[8]),
    .d(al_1315ed94[6]),
    .e(al_1315ed94[7]),
    .f(al_1315ed94[8]),
    .o(al_a24ece81));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(F@D)*~(E@C))"),
    .INIT(64'h8000080000800008))
    al_73feb8e9 (
    .a(al_a24ece81),
    .b(al_ec383fcc),
    .c(al_11033702[9]),
    .d(al_11033702[11]),
    .e(al_1315ed94[9]),
    .f(al_1315ed94[11]),
    .o(al_ff12c8b));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_ab9443b7 (
    .a(al_11033702[0]),
    .b(al_1315ed94[0]),
    .o(al_ad33515c));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_585fab01 (
    .a(al_11033702[3]),
    .b(al_1315ed94[3]),
    .o(al_d4dcd819));
  AL_MAP_LUT6 #(
    .EQN("(~B*(~(A)*~(C)*~(D)*~(E)*~(F)+~(A)*~(C)*~(D)*E*~(F)+A*~(C)*~(D)*E*~(F)+~(A)*C*~(D)*E*~(F)+~(A)*~(C)*~(D)*~(E)*F+A*~(C)*~(D)*~(E)*F+~(A)*C*~(D)*~(E)*F+A*C*~(D)*~(E)*F+~(A)*~(C)*D*~(E)*F+~(A)*~(C)*~(D)*E*F+A*~(C)*~(D)*E*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+~(A)*~(C)*D*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F))"),
    .INIT(64'h1333013300130001))
    al_455d860e (
    .a(al_ad33515c),
    .b(al_d4dcd819),
    .c(al_11033702[1]),
    .d(al_11033702[2]),
    .e(al_1315ed94[1]),
    .f(al_1315ed94[2]),
    .o(al_d69530ee));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ce8e15d (
    .a(al_11033702[3]),
    .b(al_1315ed94[3]),
    .o(al_6c403517));
  AL_MAP_LUT6 #(
    .EQN("((~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+(~B*~A)*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'h1000f100ff10fff1))
    al_e13714e4 (
    .a(al_d69530ee),
    .b(al_6c403517),
    .c(al_11033702[4]),
    .d(al_11033702[5]),
    .e(al_1315ed94[4]),
    .f(al_1315ed94[5]),
    .o(al_754ea4fe));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*(C*~A)*~(D)+~(B)*~((C*~A))*D+~(B)*(C*~A)*D+B*(C*~A)*D)"),
    .INIT(16'h7310))
    al_3c9345cf (
    .a(al_11033702[6]),
    .b(al_11033702[7]),
    .c(al_1315ed94[6]),
    .d(al_1315ed94[7]),
    .o(al_18e25363));
  AL_MAP_LUT6 #(
    .EQN("(B*(A*~(C)*~(D)*~(E)*~(F)+~(A)*~(C)*~(D)*E*~(F)+A*~(C)*~(D)*E*~(F)+A*C*~(D)*E*~(F)+~(A)*~(C)*~(D)*~(E)*F+A*~(C)*~(D)*~(E)*F+~(A)*C*~(D)*~(E)*F+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+~(A)*~(C)*~(D)*E*F+A*~(C)*~(D)*E*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+~(A)*~(C)*D*E*F+A*~(C)*D*E*F+A*C*D*E*F))"),
    .INIT(64'h8ccc08cc008c0008))
    al_ceefb38e (
    .a(al_18e25363),
    .b(al_ec383fcc),
    .c(al_11033702[8]),
    .d(al_11033702[9]),
    .e(al_1315ed94[8]),
    .f(al_1315ed94[9]),
    .o(al_37bc7186));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_a077008 (
    .a(al_b2a0a3a),
    .b(al_ad38578c),
    .c(al_11033702[21]),
    .d(al_11033702[22]),
    .o(al_e110622d));
  AL_MAP_LUT6 #(
    .EQN("(C*A*((~D*~B)*~(E)*~(F)+~((~D*~B))*E*~(F)+(~D*~B)*E*~(F)+(~D*~B)*E*F))"),
    .INIT(64'h00200000a0a00020))
    al_75783880 (
    .a(al_a0f967e6),
    .b(al_37bc7186),
    .c(al_30ecd40b),
    .d(al_2105c1a),
    .e(al_11033702[11]),
    .f(al_1315ed94[11]),
    .o(al_2219a139));
  AL_MAP_LUT6 #(
    .EQN("(~D*~C*(~(B)*(E*~A)*~(F)+~(B)*~((E*~A))*F+~(B)*(E*~A)*F+B*(E*~A)*F))"),
    .INIT(64'h0007000300010000))
    al_6ac84dc0 (
    .a(al_11033702[19]),
    .b(al_11033702[20]),
    .c(al_11033702[21]),
    .d(al_11033702[22]),
    .e(al_1315ed94[19]),
    .f(al_1315ed94[20]),
    .o(al_244bf368));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_2f9194b9 (
    .a(al_244bf368),
    .b(al_11033702[23]),
    .c(al_11033702[24]),
    .d(al_11033702[25]),
    .e(al_11033702[26]),
    .o(al_cb2a582d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_5cd9affa (
    .a(al_11033702[27]),
    .b(al_11033702[28]),
    .c(al_11033702[29]),
    .d(al_11033702[30]),
    .e(al_11033702[31]),
    .f(al_11033702[32]),
    .o(al_65ae4a67));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_f0f748ad (
    .a(al_11033702[33]),
    .b(al_11033702[36]),
    .c(al_11033702[37]),
    .d(al_11033702[38]),
    .e(al_11033702[39]),
    .f(al_11033702[40]),
    .o(al_5d4ddebc));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_54ed53ed (
    .a(al_65ae4a67),
    .b(al_5d4ddebc),
    .c(al_11033702[34]),
    .d(al_11033702[35]),
    .o(al_d5e7ffcc));
  AL_MAP_LUT6 #(
    .EQN("(D*~(~F*~(A*~(B*~(E*~C)))))"),
    .INIT(64'hff00ff002a002200))
    al_dc29d0c3 (
    .a(al_3f9c0f6c),
    .b(al_2219a139),
    .c(al_754ea4fe),
    .d(al_d5e7ffcc),
    .e(al_ff12c8b),
    .f(al_cb2a582d),
    .o(al_c61b4192));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_f08e2782 (
    .a(numerator[20]),
    .b(numerator[19]),
    .c(al_563a08a7[19]),
    .o(al_a8ba9585));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_2f65652b (
    .a(al_c61b4192),
    .b(al_a8ba9585),
    .c(start),
    .d(al_1315ed94[19]),
    .e(al_248537e7[19]),
    .o(al_9bfb1470[19]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_3c9ff229 (
    .a(al_11033702[16]),
    .b(al_1315ed94[16]),
    .o(al_a93ceae5));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_1d177e08 (
    .a(al_11033702[15]),
    .b(al_1315ed94[15]),
    .o(al_f2884563));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_db832082 (
    .a(numerator[20]),
    .b(numerator[1]),
    .c(al_563a08a7[1]),
    .o(al_1f2fd634));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_e0f43cc1 (
    .a(al_c61b4192),
    .b(al_1f2fd634),
    .c(start),
    .d(al_1315ed94[1]),
    .e(al_248537e7[1]),
    .o(al_9bfb1470[1]));
  AL_MAP_LUT6 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~((F*B))*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*(F*B)*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*(F*B)*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*(F*B)*C)"),
    .INIT(64'hcfcac5c00f0a0500))
    al_e01dd5be (
    .a(al_c61b4192),
    .b(numerator[20]),
    .c(start),
    .d(al_1315ed94[20]),
    .e(al_248537e7[20]),
    .f(al_563a08a7[20]),
    .o(al_9bfb1470[20]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_3e04c0e7 (
    .a(numerator[20]),
    .b(numerator[2]),
    .c(al_563a08a7[2]),
    .o(al_2666c71d));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_ec1b4fb9 (
    .a(al_c61b4192),
    .b(al_2666c71d),
    .c(start),
    .d(al_1315ed94[2]),
    .e(al_248537e7[2]),
    .o(al_9bfb1470[2]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_b86e3fac (
    .a(numerator[20]),
    .b(numerator[3]),
    .c(al_563a08a7[3]),
    .o(al_e662d6df));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_2ebca82 (
    .a(al_c61b4192),
    .b(al_e662d6df),
    .c(start),
    .d(al_1315ed94[3]),
    .e(al_248537e7[3]),
    .o(al_9bfb1470[3]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_1f499def (
    .a(numerator[20]),
    .b(numerator[4]),
    .c(al_563a08a7[4]),
    .o(al_c0ec79fe));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_f2e9961a (
    .a(al_c61b4192),
    .b(al_c0ec79fe),
    .c(start),
    .d(al_1315ed94[4]),
    .e(al_248537e7[4]),
    .o(al_9bfb1470[4]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_8f1711f3 (
    .a(numerator[20]),
    .b(numerator[5]),
    .c(al_563a08a7[5]),
    .o(al_91f93bf1));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_34eb6404 (
    .a(al_c61b4192),
    .b(al_91f93bf1),
    .c(start),
    .d(al_1315ed94[5]),
    .e(al_248537e7[5]),
    .o(al_9bfb1470[5]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_6e1c653d (
    .a(numerator[20]),
    .b(numerator[6]),
    .c(al_563a08a7[6]),
    .o(al_3827637d));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_dd4a87d1 (
    .a(al_c61b4192),
    .b(al_3827637d),
    .c(start),
    .d(al_1315ed94[6]),
    .e(al_248537e7[6]),
    .o(al_9bfb1470[6]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_b46e3fd7 (
    .a(numerator[20]),
    .b(numerator[7]),
    .c(al_563a08a7[7]),
    .o(al_e18beeda));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_24a1206 (
    .a(al_c61b4192),
    .b(al_e18beeda),
    .c(start),
    .d(al_1315ed94[7]),
    .e(al_248537e7[7]),
    .o(al_9bfb1470[7]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_d21f8608 (
    .a(numerator[20]),
    .b(numerator[8]),
    .c(al_563a08a7[8]),
    .o(al_c8377ec7));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_99779fac (
    .a(al_c61b4192),
    .b(al_c8377ec7),
    .c(start),
    .d(al_1315ed94[8]),
    .e(al_248537e7[8]),
    .o(al_9bfb1470[8]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_42e41119 (
    .a(numerator[20]),
    .b(numerator[9]),
    .c(al_563a08a7[9]),
    .o(al_60559583));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~(~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'h3f3a3530))
    al_1aa42175 (
    .a(al_c61b4192),
    .b(al_60559583),
    .c(start),
    .d(al_1315ed94[9]),
    .e(al_248537e7[9]),
    .o(al_9bfb1470[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b4f9e9c3 (
    .a(al_f1a38dd5),
    .b(al_327525b3[10]),
    .c(al_80e06344[10]),
    .o(al_dd9da09a[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_603d02b3 (
    .a(al_f1a38dd5),
    .b(al_327525b3[11]),
    .c(al_80e06344[11]),
    .o(al_dd9da09a[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1b69344e (
    .a(al_f1a38dd5),
    .b(al_327525b3[12]),
    .c(al_80e06344[12]),
    .o(al_dd9da09a[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6b999f16 (
    .a(al_f1a38dd5),
    .b(al_327525b3[13]),
    .c(al_80e06344[13]),
    .o(al_dd9da09a[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_37d5aed4 (
    .a(al_f1a38dd5),
    .b(al_327525b3[14]),
    .c(al_80e06344[14]),
    .o(al_dd9da09a[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1566204d (
    .a(al_f1a38dd5),
    .b(al_327525b3[15]),
    .c(al_80e06344[15]),
    .o(al_dd9da09a[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bb0704e (
    .a(al_f1a38dd5),
    .b(al_327525b3[16]),
    .c(al_80e06344[16]),
    .o(al_dd9da09a[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_918cd26d (
    .a(al_f1a38dd5),
    .b(al_327525b3[17]),
    .c(al_80e06344[17]),
    .o(al_dd9da09a[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_57add5b8 (
    .a(al_f1a38dd5),
    .b(al_327525b3[18]),
    .c(al_80e06344[18]),
    .o(al_dd9da09a[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d7e25f77 (
    .a(al_f1a38dd5),
    .b(al_327525b3[19]),
    .c(al_80e06344[19]),
    .o(al_dd9da09a[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_44e8b792 (
    .a(al_f1a38dd5),
    .b(al_327525b3[1]),
    .c(al_80e06344[1]),
    .o(al_dd9da09a[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_94078cde (
    .a(al_f1a38dd5),
    .b(al_327525b3[20]),
    .c(al_80e06344[20]),
    .o(al_dd9da09a[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c84024bf (
    .a(al_f1a38dd5),
    .b(al_327525b3[2]),
    .c(al_80e06344[2]),
    .o(al_dd9da09a[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3af7bdd7 (
    .a(al_f1a38dd5),
    .b(al_327525b3[3]),
    .c(al_80e06344[3]),
    .o(al_dd9da09a[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b9fd2bef (
    .a(al_f1a38dd5),
    .b(al_327525b3[4]),
    .c(al_80e06344[4]),
    .o(al_dd9da09a[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_99cc872 (
    .a(al_f1a38dd5),
    .b(al_327525b3[5]),
    .c(al_80e06344[5]),
    .o(al_dd9da09a[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_829c404f (
    .a(al_f1a38dd5),
    .b(al_327525b3[6]),
    .c(al_80e06344[6]),
    .o(al_dd9da09a[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a291c151 (
    .a(al_f1a38dd5),
    .b(al_327525b3[7]),
    .c(al_80e06344[7]),
    .o(al_dd9da09a[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fb2c306a (
    .a(al_f1a38dd5),
    .b(al_327525b3[8]),
    .c(al_80e06344[8]),
    .o(al_dd9da09a[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bc50cc28 (
    .a(al_f1a38dd5),
    .b(al_327525b3[9]),
    .c(al_80e06344[9]),
    .o(al_dd9da09a[9]));
  AL_DFF_0 al_3b47d798 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_55b210dc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1a38dd5));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_cf448d0 (
    .a(numerator[20]),
    .b(start),
    .c(al_f1a38dd5),
    .o(al_55b210dc));
  AL_DFF_0 al_b26d62bf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[0]));
  AL_DFF_0 al_809f7104 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[1]));
  AL_DFF_0 al_c1468025 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[2]));
  AL_DFF_0 al_c19d8344 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[3]));
  AL_DFF_0 al_ca1eda73 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[4]));
  AL_DFF_0 al_b40e8e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[8]));
  AL_DFF_0 al_2259e8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[9]));
  AL_DFF_0 al_5f624aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[10]));
  AL_DFF_0 al_d532b054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[11]));
  AL_DFF_0 al_9d987fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[12]));
  AL_DFF_0 al_220744cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[13]));
  AL_DFF_0 al_e241f44a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[14]));
  AL_DFF_0 al_897da5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[15]));
  AL_DFF_0 al_9e863954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[16]));
  AL_DFF_0 al_a186fcad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[17]));
  AL_DFF_0 al_fd544ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[0]));
  AL_DFF_0 al_21ba363c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[18]));
  AL_DFF_0 al_c602bc36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[19]));
  AL_DFF_0 al_be443a52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[20]));
  AL_DFF_0 al_961a8bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[21]));
  AL_DFF_0 al_6d594c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[22]));
  AL_DFF_0 al_5e95843a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[23]));
  AL_DFF_0 al_d701a9b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[24]));
  AL_DFF_0 al_420d26fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[25]));
  AL_DFF_0 al_eb274ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[26]));
  AL_DFF_0 al_59566ddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[27]));
  AL_DFF_0 al_40ebe0d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[1]));
  AL_DFF_0 al_88ac72e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[28]));
  AL_DFF_0 al_415d213a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[29]));
  AL_DFF_0 al_2589b38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[30]));
  AL_DFF_0 al_d3625316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[31]));
  AL_DFF_0 al_a773e9fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[32]));
  AL_DFF_0 al_b5a98930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[33]));
  AL_DFF_0 al_84e187a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[34]));
  AL_DFF_0 al_f3095820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[35]));
  AL_DFF_0 al_9b82a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[36]));
  AL_DFF_0 al_e2ab1094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[37]));
  AL_DFF_0 al_b4cd3408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[2]));
  AL_DFF_0 al_a247c67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[38]));
  AL_DFF_0 al_538bab61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[39]));
  AL_DFF_0 al_39eff7a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[20]),
    .en(1'b1),
    .sr(~start),
    .ss(1'b0),
    .q(al_11033702[40]));
  AL_DFF_0 al_16607eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[3]));
  AL_DFF_0 al_2e1082f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[4]));
  AL_DFF_0 al_806f02ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[5]));
  AL_DFF_0 al_e97bb64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[6]));
  AL_DFF_0 al_f7f2da08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[7]));
  AL_DFF_0 al_596b0fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[8]));
  AL_DFF_0 al_5cfa2c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[9]));
  AL_DFF_0 al_c56c02f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[10]));
  AL_DFF_0 al_60ec2662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[11]));
  AL_DFF_0 al_ea3f598e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[12]));
  AL_DFF_0 al_dd4ae85d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[13]));
  AL_DFF_0 al_e2aa8055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[14]));
  AL_DFF_0 al_82aa8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[15]));
  AL_DFF_0 al_7f911c70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[16]));
  AL_DFF_0 al_8908ba38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[17]));
  AL_DFF_0 al_16ad90bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[0]));
  AL_DFF_0 al_2149b062 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[18]));
  AL_DFF_0 al_56d82898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[19]));
  AL_DFF_0 al_c8bec57f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[20]));
  AL_DFF_0 al_e1044ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[1]));
  AL_DFF_0 al_16da6de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[2]));
  AL_DFF_0 al_e819e904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[3]));
  AL_DFF_0 al_4990808d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[4]));
  AL_DFF_0 al_d51e17ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[5]));
  AL_DFF_0 al_b67f884b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[6]));
  AL_DFF_0 al_ff3308ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[7]));
  AL_DFF_0 al_c1e3ea45 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[8]));
  AL_DFF_0 al_b7aa029f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[9]));
  AL_DFF_0 al_2f4f18cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[10]));
  AL_DFF_0 al_42a7eb97 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[11]));
  AL_DFF_0 al_f77c099a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[12]));
  AL_DFF_0 al_6893ba8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[13]));
  AL_DFF_0 al_d6d1e991 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[14]));
  AL_DFF_0 al_4d3bf6cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[15]));
  AL_DFF_0 al_aa8c310 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[16]));
  AL_DFF_0 al_d8095998 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[17]));
  AL_DFF_0 al_53efe64b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[0]));
  AL_DFF_0 al_68082bd4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[18]));
  AL_DFF_0 al_d9e8ef9f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[19]));
  AL_DFF_0 al_39169fb8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[20]));
  AL_DFF_0 al_26890f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[1]));
  AL_DFF_0 al_802c7023 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[2]));
  AL_DFF_0 al_9c45670 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[3]));
  AL_DFF_0 al_b0a0e999 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[4]));
  AL_DFF_0 al_739d9f2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[5]));
  AL_DFF_0 al_7f9eee7d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[6]));
  AL_DFF_0 al_741313a7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dd9da09a[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[7]));
  AL_DFF_0 al_ce6e5997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[8]));
  AL_DFF_0 al_7c322425 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[9]));
  AL_DFF_0 al_1f65ec13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[10]));
  AL_DFF_0 al_63457b5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[11]));
  AL_DFF_0 al_11fe6cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[12]));
  AL_DFF_0 al_9cfb6f54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[13]));
  AL_DFF_0 al_40b705d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[14]));
  AL_DFF_0 al_cbb21b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[15]));
  AL_DFF_0 al_a743530c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[16]));
  AL_DFF_0 al_50032887 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[17]));
  AL_DFF_0 al_5e904a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c61b4192),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[0]));
  AL_DFF_0 al_db3b2b53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[18]));
  AL_DFF_0 al_4496adb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[19]));
  AL_DFF_0 al_db38e2c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[20]));
  AL_DFF_0 al_116f1db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[1]));
  AL_DFF_0 al_6c993e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[2]));
  AL_DFF_0 al_23963ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[3]));
  AL_DFF_0 al_6c25cf29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[4]));
  AL_DFF_0 al_e7cc423c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[5]));
  AL_DFF_0 al_2c6ea385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[6]));
  AL_DFF_0 al_a356779f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[7]));
  AL_DFF_0 al_f27b108d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[8]));
  AL_DFF_0 al_d1a67c2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[9]));
  AL_DFF_0 al_a7f95d18 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[10]));
  AL_DFF_0 al_da9c9cea (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[11]));
  AL_DFF_0 al_40fd9462 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[12]));
  AL_DFF_0 al_ac95b5a9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[13]));
  AL_DFF_0 al_1a9bbf3f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[14]));
  AL_DFF_0 al_66512653 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[15]));
  AL_DFF_0 al_ec92959e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[16]));
  AL_DFF_0 al_efe05263 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[17]));
  AL_DFF_0 al_cbbb4490 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[0]));
  AL_DFF_0 al_79481707 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[18]));
  AL_DFF_0 al_ed94bd54 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[19]));
  AL_DFF_0 al_a15c98bd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[20]));
  AL_DFF_0 al_30153836 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[1]));
  AL_DFF_0 al_37ead40d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[2]));
  AL_DFF_0 al_7625712c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[3]));
  AL_DFF_0 al_2531de5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[4]));
  AL_DFF_0 al_2ccbdc6d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[5]));
  AL_DFF_0 al_2c62c395 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[6]));
  AL_DFF_0 al_ee1990ef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_50fbc01b[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_e9d64c7 (
    .a(al_1315ed94[10]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[10]),
    .o(al_50fbc01b[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_cbc5bbb8 (
    .a(al_1315ed94[11]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[11]),
    .o(al_50fbc01b[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_388f20e6 (
    .a(al_1315ed94[12]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[12]),
    .o(al_50fbc01b[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_f75a707f (
    .a(al_1315ed94[13]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[13]),
    .o(al_50fbc01b[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_20e33472 (
    .a(al_1315ed94[14]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[14]),
    .o(al_50fbc01b[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_6c3077e6 (
    .a(al_1315ed94[15]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[15]),
    .o(al_50fbc01b[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_a1004e93 (
    .a(al_1315ed94[16]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[16]),
    .o(al_50fbc01b[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_59add51 (
    .a(al_1315ed94[17]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[17]),
    .o(al_50fbc01b[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_91914bf3 (
    .a(al_1315ed94[18]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[18]),
    .o(al_50fbc01b[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_327b16fb (
    .a(al_1315ed94[19]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[19]),
    .o(al_50fbc01b[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_c45afe8c (
    .a(al_1315ed94[1]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[1]),
    .o(al_50fbc01b[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_1613fb8c (
    .a(al_1315ed94[20]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[20]),
    .o(al_50fbc01b[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_3ae6bdd1 (
    .a(al_1315ed94[2]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[2]),
    .o(al_50fbc01b[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_24a5858 (
    .a(al_1315ed94[3]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[3]),
    .o(al_50fbc01b[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_78d16bf3 (
    .a(al_1315ed94[4]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[4]),
    .o(al_50fbc01b[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_ece4c68a (
    .a(al_1315ed94[5]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[5]),
    .o(al_50fbc01b[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_a85824e4 (
    .a(al_1315ed94[6]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[6]),
    .o(al_50fbc01b[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_f3af1371 (
    .a(al_1315ed94[7]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[7]),
    .o(al_50fbc01b[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_9fe74d01 (
    .a(al_1315ed94[8]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[8]),
    .o(al_50fbc01b[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_d3702d2 (
    .a(al_1315ed94[9]),
    .b(al_4ad78cf7),
    .c(al_6e5e4cef[9]),
    .o(al_50fbc01b[9]));
  AL_DFF_0 al_4560ed77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4ad78cf7));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_1315ed94[7]),
    .b(al_11033702[7]),
    .c(al_d16993ed),
    .o({al_ae0a6293,al_248537e7[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_1315ed94[8]),
    .b(al_11033702[8]),
    .c(al_ae0a6293),
    .o({al_d07a623a,al_248537e7[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_1315ed94[9]),
    .b(al_11033702[9]),
    .c(al_d07a623a),
    .o({al_126bbf82,al_248537e7[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_1315ed94[10]),
    .b(al_11033702[10]),
    .c(al_126bbf82),
    .o({al_1aac3445,al_248537e7[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_1315ed94[11]),
    .b(al_11033702[11]),
    .c(al_1aac3445),
    .o({al_f5516224,al_248537e7[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_1315ed94[12]),
    .b(al_11033702[12]),
    .c(al_f5516224),
    .o({al_91108e0e,al_248537e7[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_1315ed94[13]),
    .b(al_11033702[13]),
    .c(al_91108e0e),
    .o({al_a4e1781b,al_248537e7[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_1315ed94[14]),
    .b(al_11033702[14]),
    .c(al_a4e1781b),
    .o({al_dc44be48,al_248537e7[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_1315ed94[15]),
    .b(al_11033702[15]),
    .c(al_dc44be48),
    .o({al_d8dd00e3,al_248537e7[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_1315ed94[16]),
    .b(al_11033702[16]),
    .c(al_d8dd00e3),
    .o({al_a0bad8f5,al_248537e7[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f5224f5b (
    .a(1'b0),
    .o({al_f39a7e9,open_n17}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_1315ed94[17]),
    .b(al_11033702[17]),
    .c(al_a0bad8f5),
    .o({al_c93e73fa,al_248537e7[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bbcbdbe (
    .a(al_1315ed94[18]),
    .b(al_11033702[18]),
    .c(al_c93e73fa),
    .o({al_6ea85cef,al_248537e7[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_216ec453 (
    .a(al_1315ed94[19]),
    .b(al_11033702[19]),
    .c(al_6ea85cef),
    .o({al_52616de9,al_248537e7[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c943a4d2 (
    .a(al_1315ed94[20]),
    .b(al_11033702[20]),
    .c(al_52616de9),
    .o({open_n18,al_248537e7[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6e3dfcf (
    .a(al_1315ed94[0]),
    .b(al_11033702[0]),
    .c(al_f39a7e9),
    .o({al_9762a925,al_248537e7[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68abff86 (
    .a(al_1315ed94[1]),
    .b(al_11033702[1]),
    .c(al_9762a925),
    .o({al_ef2ad0c3,al_248537e7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_1315ed94[2]),
    .b(al_11033702[2]),
    .c(al_ef2ad0c3),
    .o({al_e7f7dbb1,al_248537e7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_1315ed94[3]),
    .b(al_11033702[3]),
    .c(al_e7f7dbb1),
    .o({al_b1f223c3,al_248537e7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_1315ed94[4]),
    .b(al_11033702[4]),
    .c(al_b1f223c3),
    .o({al_e7086bfe,al_248537e7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_1315ed94[5]),
    .b(al_11033702[5]),
    .c(al_e7086bfe),
    .o({al_5e7e4908,al_248537e7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_1315ed94[6]),
    .b(al_11033702[6]),
    .c(al_5e7e4908),
    .o({al_d16993ed,al_248537e7[6]}));

endmodule 

