// Verilog netlist created by Tang Dynasty v5.6.60861
// Tue Oct 25 14:28:56 2022

`timescale 1ns / 1ps
module unsigned32_unsigned32_divider
  (
  clk,
  denominator,
  numerator,
  rst,
  start,
  done,
  quotient,
  remainder
  );

  input clk;
  input [31:0] denominator;
  input [43:0] numerator;
  input rst;
  input start;
  output done;
  output [43:0] quotient;
  output [31:0] remainder;

  parameter S_DEN = "UNSIGNED";
  parameter S_NUM = "UNSIGNED";
  parameter W_DEN = 32;
  parameter W_NUM = 44;
  // localparam W_CNT = 6;
  wire [5:0] al_1deac949;
  wire [5:0] al_d0dc52fd;
  wire [5:0] al_8105fe59;
  wire [74:0] al_11033702;
  wire [74:0] al_1c1b24e7;
  wire [43:0] al_1315ed94;
  wire [43:0] al_9bfb1470;
  wire [74:0] al_c67bebad;
  wire [43:0] al_327525b3;
  wire al_e583107e;
  wire al_944d9d4;
  wire al_f373539a;
  wire al_750066a4;
  wire al_74601237;
  wire al_9ea60d40;
  wire al_66e20fd7;
  wire al_c42610d7;
  wire al_aafcdc4e;
  wire al_2e8fa021;
  wire al_a190bdcc;
  wire al_75d460f3;
  wire al_47099ed2;
  wire al_90b83da;
  wire al_858ded8f;
  wire al_2485c0ac;
  wire al_b8f81b5;
  wire al_8e42eb56;
  wire al_4569ed18;
  wire al_b45ee106;
  wire al_d5a1b053;
  wire al_4be023c;
  wire al_6c2b8266;
  wire al_2f163c05;
  wire al_8b8c48b7;
  wire al_a2e92837;
  wire al_f656725a;
  wire al_28354a20;
  wire al_23e4bcdc;
  wire al_45f4f2c6;
  wire al_ddde0c42;
  wire al_6fbb2d82;
  wire al_a9d932ce;
  wire al_ecfcb3a4;
  wire al_a3626bfc;
  wire al_9031f908;
  wire al_94ad97ab;
  wire al_a6a5fe68;
  wire al_467db6bc;
  wire al_2c4eadf4;
  wire al_136010db;
  wire al_3e351de0;
  wire al_89cd14a1;
  wire al_7e7ca026;
  wire al_cde0b283;
  wire al_114eba31;
  wire al_c61b4192;
  wire al_2ea6dadb;
  wire al_3ceb5ea8;
  wire al_48b4b189;
  wire al_698e288c;
  wire al_6e8802d0;
  wire al_4ebc85a1;
  wire al_64605a2;
  wire al_77d55c19;
  wire al_5ff7b23c;
  wire al_55fd905a;
  wire al_db8535a1;
  wire al_6a8a512a;
  wire al_2cd2cfbe;
  wire al_143f80fc;
  wire al_d2146a53;
  wire al_f2f5c5f9;
  wire al_9f41e076;
  wire al_a7e41d98;
  wire al_7840e15b;
  wire al_7a9fa9c2;
  wire al_4996a689;
  wire al_66690ee5;
  wire al_f0f82df9;
  wire al_b902623;
  wire al_cbd50f66;
  wire al_e50371ba;
  wire al_6e8630b9;
  wire al_7556f838;
  wire al_2d9bc500;
  wire al_90cd446f;
  wire al_7cc72b1c;
  wire al_a81bbf88;
  wire al_7e75500b;
  wire al_f0003727;
  wire al_70feb7d0;
  wire al_7b6e6516;
  wire al_dfe291fa;
  wire al_600a9d2d;
  wire al_ba48675f;
  wire al_65a3cdd3;
  wire al_a254748;
  wire al_df3a8195;
  wire al_3e41d67f;
  wire al_9f1c02e3;
  wire al_b720b7ea;
  wire al_76496599;
  wire al_c9ed4023;
  wire al_ee6f5055;
  wire al_3125689a;
  wire al_2d31db3e;
  wire al_83a87c3b;
  wire al_ffe16699;
  wire al_f00f5cc4;
  wire al_2d062697;
  wire al_e84dfba;
  wire al_daac6179;
  wire al_b6bcb7c8;

  AL_MAP_LUT6 #(
    .EQN("(~A*~(~F*~E*~D*~C*~B))"),
    .INIT(64'h5555555555555554))
    al_f17cd423 (
    .a(al_1deac949[0]),
    .b(al_1deac949[1]),
    .c(al_1deac949[2]),
    .d(al_1deac949[3]),
    .e(al_1deac949[4]),
    .f(al_1deac949[5]),
    .o(al_8105fe59[0]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_b5f6bee4 (
    .a(al_8105fe59[0]),
    .b(start),
    .o(al_d0dc52fd[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    al_147e6a1b (
    .a(al_3ceb5ea8),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .o(al_d0dc52fd[1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(C*B)))"),
    .INIT(16'h2a80))
    al_c8620855 (
    .a(al_3ceb5ea8),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .o(al_d0dc52fd[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_6614de08 (
    .a(al_2ea6dadb),
    .b(al_1deac949[1]),
    .c(al_1deac949[4]),
    .d(al_1deac949[5]),
    .o(al_114eba31));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_2c5ab42c (
    .a(al_114eba31),
    .b(start),
    .o(al_3ceb5ea8));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@(D*C*B)))"),
    .INIT(32'h2aaa8000))
    al_ae122613 (
    .a(al_3ceb5ea8),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .e(al_1deac949[3]),
    .o(al_d0dc52fd[3]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_6dc5f615 (
    .a(al_2ea6dadb),
    .b(start),
    .c(al_1deac949[1]),
    .d(al_1deac949[4]),
    .o(al_d0dc52fd[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_79196817 (
    .a(al_1deac949[0]),
    .b(al_1deac949[2]),
    .c(al_1deac949[3]),
    .o(al_2ea6dadb));
  AL_MAP_LUT5 #(
    .EQN("(~B*(A*C*D*~(E)+~(A)*~(C)*~(D)*E+~(A)*C*~(D)*E+A*C*~(D)*E+~(A)*~(C)*D*E+A*~(C)*D*E+~(A)*C*D*E))"),
    .INIT(32'h13312000))
    al_e3df142c (
    .a(al_2ea6dadb),
    .b(start),
    .c(al_1deac949[1]),
    .d(al_1deac949[4]),
    .e(al_1deac949[5]),
    .o(al_d0dc52fd[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7885a4da (
    .a(denominator[0]),
    .b(start),
    .c(al_11033702[44]),
    .o(al_1c1b24e7[43]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_d4d1b5a8 (
    .a(denominator[1]),
    .b(start),
    .c(al_11033702[45]),
    .o(al_1c1b24e7[44]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8180372b (
    .a(denominator[2]),
    .b(start),
    .c(al_11033702[46]),
    .o(al_1c1b24e7[45]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f5c2596c (
    .a(denominator[3]),
    .b(start),
    .c(al_11033702[47]),
    .o(al_1c1b24e7[46]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_21badd87 (
    .a(denominator[4]),
    .b(start),
    .c(al_11033702[48]),
    .o(al_1c1b24e7[47]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1f53bb72 (
    .a(denominator[5]),
    .b(start),
    .c(al_11033702[49]),
    .o(al_1c1b24e7[48]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b0febaf3 (
    .a(denominator[6]),
    .b(start),
    .c(al_11033702[50]),
    .o(al_1c1b24e7[49]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1278d55d (
    .a(denominator[7]),
    .b(start),
    .c(al_11033702[51]),
    .o(al_1c1b24e7[50]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_edab9316 (
    .a(denominator[8]),
    .b(start),
    .c(al_11033702[52]),
    .o(al_1c1b24e7[51]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1732f7be (
    .a(denominator[9]),
    .b(start),
    .c(al_11033702[53]),
    .o(al_1c1b24e7[52]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a0c3193 (
    .a(denominator[10]),
    .b(start),
    .c(al_11033702[54]),
    .o(al_1c1b24e7[53]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7ac48cbe (
    .a(denominator[11]),
    .b(start),
    .c(al_11033702[55]),
    .o(al_1c1b24e7[54]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1580b4d7 (
    .a(denominator[12]),
    .b(start),
    .c(al_11033702[56]),
    .o(al_1c1b24e7[55]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b676dfb6 (
    .a(denominator[13]),
    .b(start),
    .c(al_11033702[57]),
    .o(al_1c1b24e7[56]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a1d1fbd0 (
    .a(denominator[14]),
    .b(start),
    .c(al_11033702[58]),
    .o(al_1c1b24e7[57]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_95aaa47a (
    .a(denominator[15]),
    .b(start),
    .c(al_11033702[59]),
    .o(al_1c1b24e7[58]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1eec55a5 (
    .a(denominator[16]),
    .b(start),
    .c(al_11033702[60]),
    .o(al_1c1b24e7[59]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8c58688c (
    .a(denominator[17]),
    .b(start),
    .c(al_11033702[61]),
    .o(al_1c1b24e7[60]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_99dd0529 (
    .a(denominator[18]),
    .b(start),
    .c(al_11033702[62]),
    .o(al_1c1b24e7[61]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_fed56650 (
    .a(denominator[19]),
    .b(start),
    .c(al_11033702[63]),
    .o(al_1c1b24e7[62]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_cb5602ba (
    .a(denominator[20]),
    .b(start),
    .c(al_11033702[64]),
    .o(al_1c1b24e7[63]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_864b0d81 (
    .a(denominator[21]),
    .b(start),
    .c(al_11033702[65]),
    .o(al_1c1b24e7[64]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a785325 (
    .a(denominator[22]),
    .b(start),
    .c(al_11033702[66]),
    .o(al_1c1b24e7[65]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_3208aa3 (
    .a(denominator[23]),
    .b(start),
    .c(al_11033702[67]),
    .o(al_1c1b24e7[66]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_538719ae (
    .a(denominator[24]),
    .b(start),
    .c(al_11033702[68]),
    .o(al_1c1b24e7[67]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f420e917 (
    .a(denominator[25]),
    .b(start),
    .c(al_11033702[69]),
    .o(al_1c1b24e7[68]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_97af0053 (
    .a(denominator[26]),
    .b(start),
    .c(al_11033702[70]),
    .o(al_1c1b24e7[69]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_169c3164 (
    .a(denominator[27]),
    .b(start),
    .c(al_11033702[71]),
    .o(al_1c1b24e7[70]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_890551f8 (
    .a(denominator[28]),
    .b(start),
    .c(al_11033702[72]),
    .o(al_1c1b24e7[71]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_ba401912 (
    .a(denominator[29]),
    .b(start),
    .c(al_11033702[73]),
    .o(al_1c1b24e7[72]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_39a194b8 (
    .a(denominator[30]),
    .b(start),
    .c(al_11033702[74]),
    .o(al_1c1b24e7[73]));
  AL_DFF_0 al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_114eba31),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_affc23c8 (
    .a(al_c61b4192),
    .b(numerator[0]),
    .c(start),
    .d(al_1315ed94[0]),
    .e(al_c67bebad[0]),
    .o(al_9bfb1470[0]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_7e4247d5 (
    .a(al_c61b4192),
    .b(numerator[10]),
    .c(start),
    .d(al_1315ed94[10]),
    .e(al_c67bebad[10]),
    .o(al_9bfb1470[10]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_8f76e334 (
    .a(al_c61b4192),
    .b(numerator[11]),
    .c(start),
    .d(al_1315ed94[11]),
    .e(al_c67bebad[11]),
    .o(al_9bfb1470[11]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_43c29c9e (
    .a(al_c61b4192),
    .b(numerator[12]),
    .c(start),
    .d(al_1315ed94[12]),
    .e(al_c67bebad[12]),
    .o(al_9bfb1470[12]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_dcb75b0 (
    .a(al_c61b4192),
    .b(numerator[13]),
    .c(start),
    .d(al_1315ed94[13]),
    .e(al_c67bebad[13]),
    .o(al_9bfb1470[13]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_e1773c9b (
    .a(al_c61b4192),
    .b(numerator[14]),
    .c(start),
    .d(al_1315ed94[14]),
    .e(al_c67bebad[14]),
    .o(al_9bfb1470[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_8e3693cb (
    .a(al_c61b4192),
    .b(numerator[15]),
    .c(start),
    .d(al_1315ed94[15]),
    .e(al_c67bebad[15]),
    .o(al_9bfb1470[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_79948be9 (
    .a(al_c61b4192),
    .b(numerator[16]),
    .c(start),
    .d(al_1315ed94[16]),
    .e(al_c67bebad[16]),
    .o(al_9bfb1470[16]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_cd0015f2 (
    .a(al_c61b4192),
    .b(numerator[17]),
    .c(start),
    .d(al_1315ed94[17]),
    .e(al_c67bebad[17]),
    .o(al_9bfb1470[17]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_5eba52cf (
    .a(al_c61b4192),
    .b(numerator[18]),
    .c(start),
    .d(al_1315ed94[18]),
    .e(al_c67bebad[18]),
    .o(al_9bfb1470[18]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_fd435063 (
    .a(al_c61b4192),
    .b(numerator[19]),
    .c(start),
    .d(al_1315ed94[19]),
    .e(al_c67bebad[19]),
    .o(al_9bfb1470[19]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_db832082 (
    .a(al_c61b4192),
    .b(numerator[1]),
    .c(start),
    .d(al_1315ed94[1]),
    .e(al_c67bebad[1]),
    .o(al_9bfb1470[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_e01dd5be (
    .a(al_c61b4192),
    .b(numerator[20]),
    .c(start),
    .d(al_1315ed94[20]),
    .e(al_c67bebad[20]),
    .o(al_9bfb1470[20]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_3caca9c9 (
    .a(al_c61b4192),
    .b(numerator[21]),
    .c(start),
    .d(al_1315ed94[21]),
    .e(al_c67bebad[21]),
    .o(al_9bfb1470[21]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_daadae89 (
    .a(al_c61b4192),
    .b(numerator[22]),
    .c(start),
    .d(al_1315ed94[22]),
    .e(al_c67bebad[22]),
    .o(al_9bfb1470[22]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_29e14add (
    .a(al_c61b4192),
    .b(numerator[23]),
    .c(start),
    .d(al_1315ed94[23]),
    .e(al_c67bebad[23]),
    .o(al_9bfb1470[23]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_144036ec (
    .a(al_c61b4192),
    .b(numerator[24]),
    .c(start),
    .d(al_1315ed94[24]),
    .e(al_c67bebad[24]),
    .o(al_9bfb1470[24]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_b86a6dbf (
    .a(al_c61b4192),
    .b(numerator[25]),
    .c(start),
    .d(al_1315ed94[25]),
    .e(al_c67bebad[25]),
    .o(al_9bfb1470[25]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_47ac1c09 (
    .a(al_c61b4192),
    .b(numerator[26]),
    .c(start),
    .d(al_1315ed94[26]),
    .e(al_c67bebad[26]),
    .o(al_9bfb1470[26]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_248ff2e3 (
    .a(al_c61b4192),
    .b(numerator[27]),
    .c(start),
    .d(al_1315ed94[27]),
    .e(al_c67bebad[27]),
    .o(al_9bfb1470[27]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_f01911bd (
    .a(al_c61b4192),
    .b(numerator[28]),
    .c(start),
    .d(al_1315ed94[28]),
    .e(al_c67bebad[28]),
    .o(al_9bfb1470[28]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_67954d07 (
    .a(al_c61b4192),
    .b(numerator[29]),
    .c(start),
    .d(al_1315ed94[29]),
    .e(al_c67bebad[29]),
    .o(al_9bfb1470[29]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_3e04c0e7 (
    .a(al_c61b4192),
    .b(numerator[2]),
    .c(start),
    .d(al_1315ed94[2]),
    .e(al_c67bebad[2]),
    .o(al_9bfb1470[2]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_3cf932bd (
    .a(al_c61b4192),
    .b(numerator[30]),
    .c(start),
    .d(al_1315ed94[30]),
    .e(al_c67bebad[30]),
    .o(al_9bfb1470[30]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_4e4f5c0d (
    .a(al_c61b4192),
    .b(numerator[31]),
    .c(start),
    .d(al_1315ed94[31]),
    .e(al_c67bebad[31]),
    .o(al_9bfb1470[31]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_2068acfa (
    .a(al_c61b4192),
    .b(numerator[32]),
    .c(start),
    .d(al_1315ed94[32]),
    .e(al_c67bebad[32]),
    .o(al_9bfb1470[32]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_b3ebb6c2 (
    .a(al_c61b4192),
    .b(numerator[33]),
    .c(start),
    .d(al_1315ed94[33]),
    .e(al_c67bebad[33]),
    .o(al_9bfb1470[33]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_4b9f6ba7 (
    .a(al_c61b4192),
    .b(numerator[34]),
    .c(start),
    .d(al_1315ed94[34]),
    .e(al_c67bebad[34]),
    .o(al_9bfb1470[34]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_a50e6b1e (
    .a(al_c61b4192),
    .b(numerator[35]),
    .c(start),
    .d(al_1315ed94[35]),
    .e(al_c67bebad[35]),
    .o(al_9bfb1470[35]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_d603efb8 (
    .a(al_c61b4192),
    .b(numerator[36]),
    .c(start),
    .d(al_1315ed94[36]),
    .e(al_c67bebad[36]),
    .o(al_9bfb1470[36]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_aa4b1285 (
    .a(al_c61b4192),
    .b(numerator[37]),
    .c(start),
    .d(al_1315ed94[37]),
    .e(al_c67bebad[37]),
    .o(al_9bfb1470[37]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_dc908fed (
    .a(al_c61b4192),
    .b(numerator[38]),
    .c(start),
    .d(al_1315ed94[38]),
    .e(al_c67bebad[38]),
    .o(al_9bfb1470[38]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_43edc8aa (
    .a(al_c61b4192),
    .b(numerator[39]),
    .c(start),
    .d(al_1315ed94[39]),
    .e(al_c67bebad[39]),
    .o(al_9bfb1470[39]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_b86e3fac (
    .a(al_c61b4192),
    .b(numerator[3]),
    .c(start),
    .d(al_1315ed94[3]),
    .e(al_c67bebad[3]),
    .o(al_9bfb1470[3]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_a9e6fc77 (
    .a(al_c61b4192),
    .b(numerator[40]),
    .c(start),
    .d(al_1315ed94[40]),
    .e(al_c67bebad[40]),
    .o(al_9bfb1470[40]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_80104e86 (
    .a(al_c61b4192),
    .b(numerator[41]),
    .c(start),
    .d(al_1315ed94[41]),
    .e(al_c67bebad[41]),
    .o(al_9bfb1470[41]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_660f5106 (
    .a(al_11033702[6]),
    .b(al_11033702[7]),
    .c(al_11033702[11]),
    .d(al_1315ed94[6]),
    .e(al_1315ed94[7]),
    .f(al_1315ed94[11]),
    .o(al_48b4b189));
  AL_MAP_LUT6 #(
    .EQN("(~B*(~(A)*~(C)*~(D)*~(E)*~(F)+~(A)*C*~(D)*~(E)*~(F)+A*C*~(D)*~(E)*~(F)+~(A)*~(C)*D*~(E)*~(F)+A*~(C)*D*~(E)*~(F)+~(A)*C*D*~(E)*~(F)+A*C*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+~(A)*~(C)*D*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*D*E*~(F)+~(A)*~(C)*D*~(E)*F+~(A)*C*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*D*E*F))"),
    .INIT(64'h1000310033103331))
    al_1cd70283 (
    .a(al_e583107e),
    .b(al_4ebc85a1),
    .c(al_11033702[2]),
    .d(al_11033702[3]),
    .e(al_1315ed94[2]),
    .f(al_1315ed94[3]),
    .o(al_64605a2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_2cefada5 (
    .a(al_11033702[62]),
    .b(al_11033702[63]),
    .c(al_11033702[64]),
    .d(al_11033702[65]),
    .e(al_11033702[66]),
    .f(al_11033702[67]),
    .o(al_ffe16699));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_41120618 (
    .a(al_11033702[56]),
    .b(al_11033702[57]),
    .c(al_11033702[58]),
    .d(al_11033702[59]),
    .e(al_11033702[60]),
    .f(al_11033702[61]),
    .o(al_f00f5cc4));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_fca0dc05 (
    .a(al_11033702[50]),
    .b(al_11033702[51]),
    .c(al_11033702[52]),
    .d(al_11033702[53]),
    .e(al_11033702[54]),
    .f(al_11033702[55]),
    .o(al_2d062697));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_bc8f96d7 (
    .a(al_11033702[46]),
    .b(al_11033702[47]),
    .c(al_11033702[48]),
    .d(al_11033702[49]),
    .e(al_11033702[74]),
    .o(al_e84dfba));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_690677be (
    .a(al_83a87c3b),
    .b(al_ffe16699),
    .c(al_f00f5cc4),
    .d(al_2d062697),
    .e(al_e84dfba),
    .o(al_daac6179));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    al_59cda085 (
    .a(al_f0003727),
    .b(al_70feb7d0),
    .c(al_7b6e6516),
    .d(al_11033702[35]),
    .e(al_1315ed94[35]),
    .o(al_b6bcb7c8));
  AL_MAP_LUT6 #(
    .EQN("(E*~(~B*~(C*~(F*D*~A))))"),
    .INIT(64'hecfc0000fcfc0000))
    al_28bd077d (
    .a(al_f0f82df9),
    .b(al_2d9bc500),
    .c(al_b720b7ea),
    .d(al_2d31db3e),
    .e(al_daac6179),
    .f(al_b6bcb7c8),
    .o(al_c61b4192));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_fbf4e3f1 (
    .a(al_c61b4192),
    .b(numerator[42]),
    .c(start),
    .d(al_1315ed94[42]),
    .e(al_c67bebad[42]),
    .o(al_9bfb1470[42]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(~(F*~D)*~(~B*~(~E*C))))"),
    .INIT(64'h22aa02aa22220202))
    al_bc4bf817 (
    .a(al_6e8802d0),
    .b(al_64605a2),
    .c(al_11033702[4]),
    .d(al_11033702[5]),
    .e(al_1315ed94[4]),
    .f(al_1315ed94[5]),
    .o(al_77d55c19));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((C*~A))*~(D)+B*~((C*~A))*~(D)+B*(C*~A)*~(D)+B*~((C*~A))*D)"),
    .INIT(16'h8cef))
    al_9cbebc89 (
    .a(al_11033702[6]),
    .b(al_11033702[7]),
    .c(al_1315ed94[6]),
    .d(al_1315ed94[7]),
    .o(al_5ff7b23c));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*C)*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    .INIT(32'h77110701))
    al_202fa688 (
    .a(al_5ff7b23c),
    .b(al_11033702[8]),
    .c(al_11033702[9]),
    .d(al_1315ed94[8]),
    .e(al_1315ed94[9]),
    .o(al_55fd905a));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d5488821 (
    .a(al_11033702[9]),
    .b(al_1315ed94[9]),
    .o(al_db8535a1));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*~(D)*E*~(F)+(~B*~A)*~(C)*~(D)*E*~(F)+~((~B*~A))*C*~(D)*E*~(F)+~((~B*~A))*~(C)*~(D)*~(E)*F+(~B*~A)*~(C)*~(D)*~(E)*F+~((~B*~A))*C*~(D)*~(E)*F+(~B*~A)*C*~(D)*~(E)*F+~((~B*~A))*~(C)*D*~(E)*F+~((~B*~A))*~(C)*~(D)*E*F+(~B*~A)*~(C)*~(D)*E*F+~((~B*~A))*C*~(D)*E*F+(~B*~A)*C*~(D)*E*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F)"),
    .INIT(64'hefff0eff00ef000e))
    al_4df93029 (
    .a(al_55fd905a),
    .b(al_db8535a1),
    .c(al_11033702[10]),
    .d(al_11033702[11]),
    .e(al_1315ed94[10]),
    .f(al_1315ed94[11]),
    .o(al_6a8a512a));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_2e807008 (
    .a(al_11033702[12]),
    .b(al_11033702[13]),
    .c(al_11033702[14]),
    .d(al_1315ed94[12]),
    .e(al_1315ed94[13]),
    .f(al_1315ed94[14]),
    .o(al_2cd2cfbe));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_3803b937 (
    .a(al_11033702[16]),
    .b(al_11033702[17]),
    .c(al_11033702[18]),
    .d(al_1315ed94[16]),
    .e(al_1315ed94[17]),
    .f(al_1315ed94[18]),
    .o(al_143f80fc));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    al_ecaf043e (
    .a(al_2cd2cfbe),
    .b(al_143f80fc),
    .c(al_11033702[15]),
    .d(al_1315ed94[15]),
    .o(al_d2146a53));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E)"),
    .INIT(32'h088cceef))
    al_d2e0fc29 (
    .a(al_11033702[13]),
    .b(al_11033702[14]),
    .c(al_1315ed94[12]),
    .d(al_1315ed94[13]),
    .e(al_1315ed94[14]),
    .o(al_f2f5c5f9));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(~C*A))"),
    .INIT(16'hc431))
    al_8ed7c2a4 (
    .a(al_11033702[5]),
    .b(al_11033702[10]),
    .c(al_1315ed94[5]),
    .d(al_1315ed94[10]),
    .o(al_698e288c));
  AL_MAP_LUT4 #(
    .EQN("(D*(~(A)*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C))"),
    .INIT(16'h7100))
    al_794af4a6 (
    .a(al_f2f5c5f9),
    .b(al_11033702[15]),
    .c(al_1315ed94[15]),
    .d(al_143f80fc),
    .o(al_9f41e076));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_ecd2ee63 (
    .a(al_11033702[23]),
    .b(al_11033702[24]),
    .c(al_11033702[25]),
    .d(al_1315ed94[23]),
    .e(al_1315ed94[24]),
    .f(al_1315ed94[25]),
    .o(al_a7e41d98));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_787aaa28 (
    .a(al_11033702[21]),
    .b(al_11033702[22]),
    .c(al_11033702[26]),
    .d(al_1315ed94[21]),
    .e(al_1315ed94[22]),
    .f(al_1315ed94[26]),
    .o(al_7840e15b));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_4b44a220 (
    .a(al_11033702[19]),
    .b(al_11033702[20]),
    .c(al_1315ed94[19]),
    .d(al_1315ed94[20]),
    .o(al_7a9fa9c2));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_b608c2f3 (
    .a(al_a7e41d98),
    .b(al_7840e15b),
    .c(al_7a9fa9c2),
    .o(al_4996a689));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((D*~A))*~(E)*~(F)+B*~(C)*~((D*~A))*~(E)*~(F)+~(B)*C*~((D*~A))*~(E)*~(F)+B*C*~((D*~A))*~(E)*~(F)+B*~(C)*(D*~A)*~(E)*~(F)+~(B)*C*(D*~A)*~(E)*~(F)+B*C*(D*~A)*~(E)*~(F)+B*~(C)*~((D*~A))*E*~(F)+~(B)*C*~((D*~A))*E*~(F)+B*C*~((D*~A))*E*~(F)+~(B)*C*(D*~A)*E*~(F)+B*C*(D*~A)*E*~(F)+~(B)*C*~((D*~A))*~(E)*F+B*C*~((D*~A))*~(E)*F+B*C*(D*~A)*~(E)*F+B*C*~((D*~A))*E*F)"),
    .INIT(64'h80c0e0f0f8fcfeff))
    al_b8e8bf81 (
    .a(al_11033702[16]),
    .b(al_11033702[17]),
    .c(al_11033702[18]),
    .d(al_1315ed94[16]),
    .e(al_1315ed94[17]),
    .f(al_1315ed94[18]),
    .o(al_66690ee5));
  AL_MAP_LUT6 #(
    .EQN("(E*~((F*~D)*~((~B*~A))*~(C)+(F*~D)*(~B*~A)*~(C)+~((F*~D))*(~B*~A)*C+(F*~D)*(~B*~A)*C))"),
    .INIT(64'hefe00000efef0000))
    al_8c36ab1e (
    .a(al_77d55c19),
    .b(al_6a8a512a),
    .c(al_d2146a53),
    .d(al_9f41e076),
    .e(al_4996a689),
    .f(al_66690ee5),
    .o(al_f0f82df9));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((C*~A))*~(D)+B*~((C*~A))*~(D)+B*(C*~A)*~(D)+B*~((C*~A))*D)"),
    .INIT(16'h8cef))
    al_a973b61c (
    .a(al_11033702[36]),
    .b(al_11033702[37]),
    .c(al_1315ed94[36]),
    .d(al_1315ed94[37]),
    .o(al_b902623));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_5b69a9ce (
    .a(al_11033702[40]),
    .b(al_1315ed94[40]),
    .o(al_cbd50f66));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*~(D)*~(E)*~(F)+~(A)*C*~(D)*~(E)*~(F)+A*C*~(D)*~(E)*~(F)+~(A)*~(C)*D*~(E)*~(F)+A*~(C)*D*~(E)*~(F)+~(A)*C*D*~(E)*~(F)+A*C*D*~(E)*~(F)+A*C*~(D)*E*~(F)+~(A)*~(C)*D*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*D*E*~(F)+A*~(C)*D*~(E)*F+~(A)*C*D*~(E)*F+A*C*D*~(E)*F+A*C*D*E*F))"),
    .INIT(64'h2000320033203332))
    al_7c2b5b2b (
    .a(al_b902623),
    .b(al_cbd50f66),
    .c(al_11033702[38]),
    .d(al_11033702[39]),
    .e(al_1315ed94[38]),
    .f(al_1315ed94[39]),
    .o(al_e50371ba));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(F@D)*~(E@C))"),
    .INIT(64'h8000080000800008))
    al_27a6a1b4 (
    .a(al_48b4b189),
    .b(al_698e288c),
    .c(al_11033702[8]),
    .d(al_11033702[9]),
    .e(al_1315ed94[8]),
    .f(al_1315ed94[9]),
    .o(al_6e8802d0));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_164a4b2f (
    .a(al_11033702[40]),
    .b(al_1315ed94[40]),
    .o(al_6e8630b9));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+~((~B*~A))*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+(~B*~A)*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*C*D*E*F)"),
    .INIT(64'he000fe00ffe0fffe))
    al_549e9dfb (
    .a(al_e50371ba),
    .b(al_6e8630b9),
    .c(al_11033702[41]),
    .d(al_11033702[42]),
    .e(al_1315ed94[41]),
    .f(al_1315ed94[42]),
    .o(al_7556f838));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(~(A)*~(B)*~(E)+~(A)*~(B)*E+A*~(B)*E+~(A)*B*E))"),
    .INIT(32'h00070001))
    al_f709e847 (
    .a(al_7556f838),
    .b(al_11033702[43]),
    .c(al_11033702[44]),
    .d(al_11033702[45]),
    .e(al_1315ed94[43]),
    .o(al_2d9bc500));
  AL_MAP_LUT6 #(
    .EQN("(~D*~C*~(F@B)*~(E@A))"),
    .INIT(64'h0008000400020001))
    al_b43a8ac2 (
    .a(al_11033702[39]),
    .b(al_11033702[43]),
    .c(al_11033702[44]),
    .d(al_11033702[45]),
    .e(al_1315ed94[39]),
    .f(al_1315ed94[43]),
    .o(al_90cd446f));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_1fff5b03 (
    .a(al_11033702[36]),
    .b(al_11033702[38]),
    .c(al_11033702[41]),
    .d(al_1315ed94[36]),
    .e(al_1315ed94[38]),
    .f(al_1315ed94[41]),
    .o(al_7cc72b1c));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_b24bed36 (
    .a(al_11033702[37]),
    .b(al_11033702[40]),
    .c(al_11033702[42]),
    .d(al_1315ed94[37]),
    .e(al_1315ed94[40]),
    .f(al_1315ed94[42]),
    .o(al_a81bbf88));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_6a86cb2a (
    .a(al_90cd446f),
    .b(al_7cc72b1c),
    .c(al_a81bbf88),
    .o(al_7e75500b));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_2fa0851e (
    .a(al_11033702[29]),
    .b(al_11033702[32]),
    .c(al_11033702[34]),
    .d(al_1315ed94[29]),
    .e(al_1315ed94[32]),
    .f(al_1315ed94[34]),
    .o(al_f0003727));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_45f455bd (
    .a(al_11033702[28]),
    .b(al_11033702[30]),
    .c(al_11033702[33]),
    .d(al_1315ed94[28]),
    .e(al_1315ed94[30]),
    .f(al_1315ed94[33]),
    .o(al_70feb7d0));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_e9e8dee3 (
    .a(al_11033702[27]),
    .b(al_11033702[31]),
    .c(al_1315ed94[27]),
    .d(al_1315ed94[31]),
    .o(al_7b6e6516));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((~C*A))*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+~(B)*(~C*A)*D)"),
    .INIT(16'hf731))
    al_3f754603 (
    .a(al_11033702[0]),
    .b(al_11033702[1]),
    .c(al_1315ed94[0]),
    .d(al_1315ed94[1]),
    .o(al_e583107e));
  AL_MAP_LUT5 #(
    .EQN("(~((C*B*A))*~(D)*~(E)+~((C*B*A))*D*~(E)+(C*B*A)*D*~(E)+~((C*B*A))*D*E)"),
    .INIT(32'h7f00ff7f))
    al_c7e51cc5 (
    .a(al_f0003727),
    .b(al_70feb7d0),
    .c(al_7b6e6516),
    .d(al_11033702[35]),
    .e(al_1315ed94[35]),
    .o(al_dfe291fa));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E)"),
    .INIT(32'h088cceef))
    al_d845b45c (
    .a(al_11033702[28]),
    .b(al_11033702[29]),
    .c(al_1315ed94[27]),
    .d(al_1315ed94[28]),
    .e(al_1315ed94[29]),
    .o(al_600a9d2d));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    al_d7146b18 (
    .a(al_11033702[31]),
    .b(al_11033702[32]),
    .c(al_1315ed94[31]),
    .d(al_1315ed94[32]),
    .o(al_ba48675f));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    al_f6b0d4f0 (
    .a(al_11033702[32]),
    .b(al_11033702[33]),
    .c(al_1315ed94[32]),
    .d(al_1315ed94[33]),
    .o(al_65a3cdd3));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_4ac30d89 (
    .a(al_11033702[31]),
    .b(al_1315ed94[31]),
    .o(al_a254748));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_5f86357c (
    .a(al_11033702[4]),
    .b(al_1315ed94[4]),
    .o(al_4ebc85a1));
  AL_MAP_LUT6 #(
    .EQN("(C*~(B*~(~D*(~(A)*~(E)*~(F)+~(A)*~(E)*F+A*~(E)*F+~(A)*E*F))))"),
    .INIT(64'h307030f030303070))
    al_df72ce56 (
    .a(al_600a9d2d),
    .b(al_ba48675f),
    .c(al_65a3cdd3),
    .d(al_a254748),
    .e(al_11033702[30]),
    .f(al_1315ed94[30]),
    .o(al_df3a8195));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    al_63002939 (
    .a(al_11033702[33]),
    .b(al_11033702[34]),
    .c(al_1315ed94[33]),
    .d(al_1315ed94[34]),
    .o(al_3e41d67f));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    al_5fde6d16 (
    .a(al_11033702[34]),
    .b(al_11033702[35]),
    .c(al_1315ed94[34]),
    .d(al_1315ed94[35]),
    .o(al_9f1c02e3));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*~(E*~(D*~C))))"),
    .INIT(32'ha2aa2222))
    al_8f4b54a (
    .a(al_7e75500b),
    .b(al_dfe291fa),
    .c(al_df3a8195),
    .d(al_3e41d67f),
    .e(al_9f1c02e3),
    .o(al_b720b7ea));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((D*~A))*~(E)*~(F)+B*~(C)*~((D*~A))*~(E)*~(F)+~(B)*C*~((D*~A))*~(E)*~(F)+B*C*~((D*~A))*~(E)*~(F)+B*~(C)*(D*~A)*~(E)*~(F)+~(B)*C*(D*~A)*~(E)*~(F)+B*C*(D*~A)*~(E)*~(F)+B*~(C)*~((D*~A))*E*~(F)+~(B)*C*~((D*~A))*E*~(F)+B*C*~((D*~A))*E*~(F)+~(B)*C*(D*~A)*E*~(F)+B*C*(D*~A)*E*~(F)+~(B)*C*~((D*~A))*~(E)*F+B*C*~((D*~A))*~(E)*F+B*C*(D*~A)*~(E)*F+B*C*~((D*~A))*E*F)"),
    .INIT(64'h80c0e0f0f8fcfeff))
    al_26f534bc (
    .a(al_11033702[19]),
    .b(al_11033702[20]),
    .c(al_11033702[21]),
    .d(al_1315ed94[19]),
    .e(al_1315ed94[20]),
    .f(al_1315ed94[21]),
    .o(al_76496599));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    al_99ea4847 (
    .a(al_11033702[23]),
    .b(al_11033702[24]),
    .c(al_1315ed94[23]),
    .d(al_1315ed94[24]),
    .o(al_c9ed4023));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    al_62cf421b (
    .a(al_11033702[24]),
    .b(al_11033702[25]),
    .c(al_1315ed94[24]),
    .d(al_1315ed94[25]),
    .o(al_ee6f5055));
  AL_MAP_LUT6 #(
    .EQN("(C*~(B*~(F*(~(A)*~(D)*~(E)+~(A)*~(D)*E+A*~(D)*E+~(A)*D*E))))"),
    .INIT(64'h70f0307030303030))
    al_f5aa2d57 (
    .a(al_76496599),
    .b(al_c9ed4023),
    .c(al_ee6f5055),
    .d(al_11033702[22]),
    .e(al_1315ed94[22]),
    .f(al_a7e41d98),
    .o(al_3125689a));
  AL_MAP_LUT5 #(
    .EQN("(C*~((~(D*~B)*~A))*~(E)+~(C)*(~(D*~B)*~A)*~(E)+C*(~(D*~B)*~A)*~(E)+C*(~(D*~B)*~A)*E)"),
    .INIT(32'h4050f4f5))
    al_dc37d187 (
    .a(al_3125689a),
    .b(al_11033702[25]),
    .c(al_11033702[26]),
    .d(al_1315ed94[25]),
    .e(al_1315ed94[26]),
    .o(al_2d31db3e));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_dfadc297 (
    .a(al_11033702[68]),
    .b(al_11033702[69]),
    .c(al_11033702[70]),
    .d(al_11033702[71]),
    .e(al_11033702[72]),
    .f(al_11033702[73]),
    .o(al_83a87c3b));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_bafb7113 (
    .a(al_c61b4192),
    .b(numerator[43]),
    .c(start),
    .d(al_1315ed94[43]),
    .e(al_c67bebad[43]),
    .o(al_9bfb1470[43]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_1f499def (
    .a(al_c61b4192),
    .b(numerator[4]),
    .c(start),
    .d(al_1315ed94[4]),
    .e(al_c67bebad[4]),
    .o(al_9bfb1470[4]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_8f1711f3 (
    .a(al_c61b4192),
    .b(numerator[5]),
    .c(start),
    .d(al_1315ed94[5]),
    .e(al_c67bebad[5]),
    .o(al_9bfb1470[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_6e1c653d (
    .a(al_c61b4192),
    .b(numerator[6]),
    .c(start),
    .d(al_1315ed94[6]),
    .e(al_c67bebad[6]),
    .o(al_9bfb1470[6]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_b46e3fd7 (
    .a(al_c61b4192),
    .b(numerator[7]),
    .c(start),
    .d(al_1315ed94[7]),
    .e(al_c67bebad[7]),
    .o(al_9bfb1470[7]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_d21f8608 (
    .a(al_c61b4192),
    .b(numerator[8]),
    .c(start),
    .d(al_1315ed94[8]),
    .e(al_c67bebad[8]),
    .o(al_9bfb1470[8]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_42e41119 (
    .a(al_c61b4192),
    .b(numerator[9]),
    .c(start),
    .d(al_1315ed94[9]),
    .e(al_c67bebad[9]),
    .o(al_9bfb1470[9]));
  AL_DFF_0 al_b26d62bf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[0]));
  AL_DFF_0 al_809f7104 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[1]));
  AL_DFF_0 al_c1468025 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[2]));
  AL_DFF_0 al_c19d8344 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[3]));
  AL_DFF_0 al_ca1eda73 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[4]));
  AL_DFF_0 al_fa89b429 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[5]));
  AL_DFF_0 al_b40e8e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[8]));
  AL_DFF_0 al_2259e8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[9]));
  AL_DFF_0 al_5f624aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[10]));
  AL_DFF_0 al_d532b054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[11]));
  AL_DFF_0 al_9d987fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[12]));
  AL_DFF_0 al_220744cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[13]));
  AL_DFF_0 al_e241f44a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[14]));
  AL_DFF_0 al_897da5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[15]));
  AL_DFF_0 al_9e863954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[16]));
  AL_DFF_0 al_a186fcad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[17]));
  AL_DFF_0 al_fd544ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[0]));
  AL_DFF_0 al_21ba363c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[18]));
  AL_DFF_0 al_c602bc36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[19]));
  AL_DFF_0 al_be443a52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[21]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[20]));
  AL_DFF_0 al_961a8bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[22]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[21]));
  AL_DFF_0 al_6d594c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[23]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[22]));
  AL_DFF_0 al_5e95843a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[24]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[23]));
  AL_DFF_0 al_d701a9b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[25]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[24]));
  AL_DFF_0 al_420d26fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[26]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[25]));
  AL_DFF_0 al_eb274ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[27]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[26]));
  AL_DFF_0 al_59566ddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[28]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[27]));
  AL_DFF_0 al_40ebe0d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[1]));
  AL_DFF_0 al_88ac72e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[29]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[28]));
  AL_DFF_0 al_415d213a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[30]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[29]));
  AL_DFF_0 al_2589b38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[31]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[30]));
  AL_DFF_0 al_d3625316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[32]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[31]));
  AL_DFF_0 al_a773e9fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[33]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[32]));
  AL_DFF_0 al_b5a98930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[34]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[33]));
  AL_DFF_0 al_84e187a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[35]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[34]));
  AL_DFF_0 al_f3095820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[36]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[35]));
  AL_DFF_0 al_9b82a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[37]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[36]));
  AL_DFF_0 al_e2ab1094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[38]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[37]));
  AL_DFF_0 al_b4cd3408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[2]));
  AL_DFF_0 al_a247c67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[39]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[38]));
  AL_DFF_0 al_538bab61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[40]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[39]));
  AL_DFF_0 al_39eff7a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[41]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[40]));
  AL_DFF_0 al_da740eac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[42]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[41]));
  AL_DFF_0 al_a1f5e6e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[43]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[42]));
  AL_DFF_0 al_73905df6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[43]));
  AL_DFF_0 al_7587b9d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[44]));
  AL_DFF_0 al_cb0b2132 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[45]));
  AL_DFF_0 al_79136648 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[46]));
  AL_DFF_0 al_a8eb1e63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[47]));
  AL_DFF_0 al_16607eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[3]));
  AL_DFF_0 al_b20ad0fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[48]));
  AL_DFF_0 al_6b481302 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[49]));
  AL_DFF_0 al_aa48a4a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[50]));
  AL_DFF_0 al_16453eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[51]));
  AL_DFF_0 al_78700b2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[52]));
  AL_DFF_0 al_3ec4517b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[53]));
  AL_DFF_0 al_f742b91d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[54]));
  AL_DFF_0 al_63888a93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[55]));
  AL_DFF_0 al_3da78364 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[56]));
  AL_DFF_0 al_3d3489ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[57]));
  AL_DFF_0 al_2e1082f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[4]));
  AL_DFF_0 al_d5896133 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[58]));
  AL_DFF_0 al_6713d36c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[59]));
  AL_DFF_0 al_498618ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[60]));
  AL_DFF_0 al_f25bea6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[61]));
  AL_DFF_0 al_2e792170 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[62]));
  AL_DFF_0 al_10e927f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[63]));
  AL_DFF_0 al_6cdaad66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[64]));
  AL_DFF_0 al_428372bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[65]));
  AL_DFF_0 al_f8209620 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[66]));
  AL_DFF_0 al_96ae94d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[67]));
  AL_DFF_0 al_806f02ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[5]));
  AL_DFF_0 al_be0c1a24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[68]));
  AL_DFF_0 al_a5d841b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[69]));
  AL_DFF_0 al_b6808dcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[70]));
  AL_DFF_0 al_5fd20133 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[71]));
  AL_DFF_0 al_57550c35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[72]));
  AL_DFF_0 al_a08195e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[73]));
  AL_DFF_0 al_8c7f06d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[31]),
    .en(1'b1),
    .sr(~start),
    .ss(1'b0),
    .q(al_11033702[74]));
  AL_DFF_0 al_e97bb64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[6]));
  AL_DFF_0 al_f7f2da08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[7]));
  AL_DFF_0 al_596b0fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[8]));
  AL_DFF_0 al_5cfa2c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[9]));
  AL_DFF_0 al_c56c02f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[10]));
  AL_DFF_0 al_60ec2662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[11]));
  AL_DFF_0 al_ea3f598e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[12]));
  AL_DFF_0 al_dd4ae85d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[13]));
  AL_DFF_0 al_e2aa8055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[14]));
  AL_DFF_0 al_82aa8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[15]));
  AL_DFF_0 al_7f911c70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[16]));
  AL_DFF_0 al_8908ba38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[17]));
  AL_DFF_0 al_16ad90bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[0]));
  AL_DFF_0 al_2149b062 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[18]));
  AL_DFF_0 al_56d82898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[19]));
  AL_DFF_0 al_c8bec57f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[20]));
  AL_DFF_0 al_1f071837 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[21]));
  AL_DFF_0 al_9acbb644 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[22]));
  AL_DFF_0 al_286bd0de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[23]));
  AL_DFF_0 al_7e8bb9f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[24]));
  AL_DFF_0 al_d4e324dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[25]));
  AL_DFF_0 al_bcaf406d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[26]));
  AL_DFF_0 al_20d194ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[27]));
  AL_DFF_0 al_e1044ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[1]));
  AL_DFF_0 al_6402198 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[28]));
  AL_DFF_0 al_3f7239b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[29]));
  AL_DFF_0 al_33cd891 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[30]));
  AL_DFF_0 al_28b9e853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[31]));
  AL_DFF_0 al_2da6eeb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[32]));
  AL_DFF_0 al_cca00973 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[33]));
  AL_DFF_0 al_6bc4a040 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[34]));
  AL_DFF_0 al_7cf6bbec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[35]));
  AL_DFF_0 al_3b3f2d26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[36]));
  AL_DFF_0 al_dc5b9d24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[37]));
  AL_DFF_0 al_16da6de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[2]));
  AL_DFF_0 al_faa19bbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[38]));
  AL_DFF_0 al_33941afe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[39]));
  AL_DFF_0 al_859d7b36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[40]));
  AL_DFF_0 al_7f8ef6ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[41]));
  AL_DFF_0 al_efcfba42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[42]));
  AL_DFF_0 al_add7811b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[43]));
  AL_DFF_0 al_e819e904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[3]));
  AL_DFF_0 al_4990808d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[4]));
  AL_DFF_0 al_d51e17ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[5]));
  AL_DFF_0 al_b67f884b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[6]));
  AL_DFF_0 al_ff3308ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[7]));
  AL_DFF_0 al_c1e3ea45 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[8]));
  AL_DFF_0 al_b7aa029f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[9]));
  AL_DFF_0 al_2f4f18cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[10]));
  AL_DFF_0 al_42a7eb97 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[11]));
  AL_DFF_0 al_f77c099a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[12]));
  AL_DFF_0 al_6893ba8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[13]));
  AL_DFF_0 al_d6d1e991 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[14]));
  AL_DFF_0 al_4d3bf6cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[15]));
  AL_DFF_0 al_aa8c310 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[16]));
  AL_DFF_0 al_d8095998 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[17]));
  AL_DFF_0 al_53efe64b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[0]));
  AL_DFF_0 al_68082bd4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[18]));
  AL_DFF_0 al_d9e8ef9f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[19]));
  AL_DFF_0 al_39169fb8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[20]));
  AL_DFF_0 al_c179532 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[21]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[21]));
  AL_DFF_0 al_7d105784 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[22]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[22]));
  AL_DFF_0 al_573a0a58 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[23]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[23]));
  AL_DFF_0 al_d0deffcb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[24]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[24]));
  AL_DFF_0 al_150254f9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[25]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[25]));
  AL_DFF_0 al_47f1ba67 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[26]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[26]));
  AL_DFF_0 al_3f6c28d5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[27]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[27]));
  AL_DFF_0 al_26890f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[1]));
  AL_DFF_0 al_930b6560 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[28]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[28]));
  AL_DFF_0 al_46a886ac (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[29]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[29]));
  AL_DFF_0 al_5c18d1b4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[30]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[30]));
  AL_DFF_0 al_f94ac09a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[31]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[31]));
  AL_DFF_0 al_4e65699f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[32]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[32]));
  AL_DFF_0 al_e18c69c7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[33]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[33]));
  AL_DFF_0 al_e1d2b0c2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[34]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[34]));
  AL_DFF_0 al_58830fc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[35]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[35]));
  AL_DFF_0 al_d9d78798 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[36]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[36]));
  AL_DFF_0 al_7013bc9a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[37]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[37]));
  AL_DFF_0 al_802c7023 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[2]));
  AL_DFF_0 al_436ca8bb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[38]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[38]));
  AL_DFF_0 al_4ccfd875 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[39]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[39]));
  AL_DFF_0 al_bb5d438b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[40]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[40]));
  AL_DFF_0 al_3f7dcd40 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[41]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[41]));
  AL_DFF_0 al_c25f43fe (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[42]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[42]));
  AL_DFF_0 al_35c2d44e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[43]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[43]));
  AL_DFF_0 al_9c45670 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[3]));
  AL_DFF_0 al_b0a0e999 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[4]));
  AL_DFF_0 al_739d9f2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[5]));
  AL_DFF_0 al_7f9eee7d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[6]));
  AL_DFF_0 al_741313a7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[7]));
  AL_DFF_0 al_ce6e5997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[8]));
  AL_DFF_0 al_7c322425 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[9]));
  AL_DFF_0 al_1f65ec13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[10]));
  AL_DFF_0 al_63457b5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[11]));
  AL_DFF_0 al_11fe6cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[12]));
  AL_DFF_0 al_9cfb6f54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[13]));
  AL_DFF_0 al_40b705d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[14]));
  AL_DFF_0 al_cbb21b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[15]));
  AL_DFF_0 al_a743530c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[16]));
  AL_DFF_0 al_50032887 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[17]));
  AL_DFF_0 al_5e904a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c61b4192),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[0]));
  AL_DFF_0 al_db3b2b53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[18]));
  AL_DFF_0 al_4496adb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[19]));
  AL_DFF_0 al_db38e2c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[20]));
  AL_DFF_0 al_b910420c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[21]));
  AL_DFF_0 al_90d7e42b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[21]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[22]));
  AL_DFF_0 al_f16a60a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[22]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[23]));
  AL_DFF_0 al_91adf23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[23]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[24]));
  AL_DFF_0 al_77ecd5d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[24]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[25]));
  AL_DFF_0 al_149f3658 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[25]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[26]));
  AL_DFF_0 al_8734a4b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[26]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[27]));
  AL_DFF_0 al_116f1db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[1]));
  AL_DFF_0 al_5bba43cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[27]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[28]));
  AL_DFF_0 al_505e168f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[28]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[29]));
  AL_DFF_0 al_a288ce99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[29]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[30]));
  AL_DFF_0 al_930333c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[30]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[31]));
  AL_DFF_0 al_5d27e954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[31]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[32]));
  AL_DFF_0 al_f0da03a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[32]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[33]));
  AL_DFF_0 al_c8a0e628 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[33]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[34]));
  AL_DFF_0 al_f689feb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[34]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[35]));
  AL_DFF_0 al_27f9e709 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[35]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[36]));
  AL_DFF_0 al_28d079d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[36]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[37]));
  AL_DFF_0 al_6c993e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[2]));
  AL_DFF_0 al_be3e1444 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[37]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[38]));
  AL_DFF_0 al_79186d83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[38]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[39]));
  AL_DFF_0 al_8a46cd85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[39]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[40]));
  AL_DFF_0 al_aa53ffe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[40]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[41]));
  AL_DFF_0 al_4203609d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[41]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[42]));
  AL_DFF_0 al_40bed0ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[42]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[43]));
  AL_DFF_0 al_23963ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[3]));
  AL_DFF_0 al_6c25cf29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[4]));
  AL_DFF_0 al_e7cc423c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[5]));
  AL_DFF_0 al_2c6ea385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[6]));
  AL_DFF_0 al_a356779f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[7]));
  AL_DFF_0 al_f27b108d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[8]));
  AL_DFF_0 al_d1a67c2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[9]));
  AL_DFF_0 al_a7f95d18 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[10]));
  AL_DFF_0 al_da9c9cea (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[11]));
  AL_DFF_0 al_40fd9462 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[12]));
  AL_DFF_0 al_ac95b5a9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[13]));
  AL_DFF_0 al_1a9bbf3f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[14]));
  AL_DFF_0 al_66512653 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[15]));
  AL_DFF_0 al_ec92959e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[16]));
  AL_DFF_0 al_efe05263 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[17]));
  AL_DFF_0 al_cbbb4490 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[0]));
  AL_DFF_0 al_79481707 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[18]));
  AL_DFF_0 al_ed94bd54 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[19]));
  AL_DFF_0 al_a15c98bd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[20]));
  AL_DFF_0 al_131a28da (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[21]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[21]));
  AL_DFF_0 al_73557a1d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[22]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[22]));
  AL_DFF_0 al_a7de7e20 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[23]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[23]));
  AL_DFF_0 al_4c32dd42 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[24]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[24]));
  AL_DFF_0 al_e05106af (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[25]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[25]));
  AL_DFF_0 al_2d9f3ce8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[26]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[26]));
  AL_DFF_0 al_de36f4d0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[27]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[27]));
  AL_DFF_0 al_30153836 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[1]));
  AL_DFF_0 al_f763c3ab (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[28]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[28]));
  AL_DFF_0 al_f3dc4f4c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[29]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[29]));
  AL_DFF_0 al_d8cfba43 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[30]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[30]));
  AL_DFF_0 al_d6316b06 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[31]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[31]));
  AL_DFF_0 al_37ead40d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[2]));
  AL_DFF_0 al_7625712c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[3]));
  AL_DFF_0 al_2531de5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[4]));
  AL_DFF_0 al_2ccbdc6d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[5]));
  AL_DFF_0 al_2c62c395 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[6]));
  AL_DFF_0 al_ee1990ef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_1315ed94[7]),
    .b(al_11033702[7]),
    .c(al_aafcdc4e),
    .o({al_2e8fa021,al_c67bebad[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_1315ed94[8]),
    .b(al_11033702[8]),
    .c(al_2e8fa021),
    .o({al_a190bdcc,al_c67bebad[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_1315ed94[9]),
    .b(al_11033702[9]),
    .c(al_a190bdcc),
    .o({al_75d460f3,al_c67bebad[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_1315ed94[10]),
    .b(al_11033702[10]),
    .c(al_75d460f3),
    .o({al_47099ed2,al_c67bebad[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_1315ed94[11]),
    .b(al_11033702[11]),
    .c(al_47099ed2),
    .o({al_90b83da,al_c67bebad[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_1315ed94[12]),
    .b(al_11033702[12]),
    .c(al_90b83da),
    .o({al_858ded8f,al_c67bebad[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_1315ed94[13]),
    .b(al_11033702[13]),
    .c(al_858ded8f),
    .o({al_2485c0ac,al_c67bebad[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_1315ed94[14]),
    .b(al_11033702[14]),
    .c(al_2485c0ac),
    .o({al_b8f81b5,al_c67bebad[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_1315ed94[15]),
    .b(al_11033702[15]),
    .c(al_b8f81b5),
    .o({al_8e42eb56,al_c67bebad[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_1315ed94[16]),
    .b(al_11033702[16]),
    .c(al_8e42eb56),
    .o({al_4569ed18,al_c67bebad[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f5224f5b (
    .a(1'b0),
    .o({al_944d9d4,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_1315ed94[17]),
    .b(al_11033702[17]),
    .c(al_4569ed18),
    .o({al_b45ee106,al_c67bebad[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bbcbdbe (
    .a(al_1315ed94[18]),
    .b(al_11033702[18]),
    .c(al_b45ee106),
    .o({al_d5a1b053,al_c67bebad[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_216ec453 (
    .a(al_1315ed94[19]),
    .b(al_11033702[19]),
    .c(al_d5a1b053),
    .o({al_4be023c,al_c67bebad[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c943a4d2 (
    .a(al_1315ed94[20]),
    .b(al_11033702[20]),
    .c(al_4be023c),
    .o({al_6c2b8266,al_c67bebad[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_920ee641 (
    .a(al_1315ed94[21]),
    .b(al_11033702[21]),
    .c(al_6c2b8266),
    .o({al_2f163c05,al_c67bebad[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e359bb16 (
    .a(al_1315ed94[22]),
    .b(al_11033702[22]),
    .c(al_2f163c05),
    .o({al_8b8c48b7,al_c67bebad[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a6af83b3 (
    .a(al_1315ed94[23]),
    .b(al_11033702[23]),
    .c(al_8b8c48b7),
    .o({al_a2e92837,al_c67bebad[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_717da7cc (
    .a(al_1315ed94[24]),
    .b(al_11033702[24]),
    .c(al_a2e92837),
    .o({al_f656725a,al_c67bebad[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_916a9569 (
    .a(al_1315ed94[25]),
    .b(al_11033702[25]),
    .c(al_f656725a),
    .o({al_28354a20,al_c67bebad[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b53f57fa (
    .a(al_1315ed94[26]),
    .b(al_11033702[26]),
    .c(al_28354a20),
    .o({al_23e4bcdc,al_c67bebad[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6e3dfcf (
    .a(al_1315ed94[0]),
    .b(al_11033702[0]),
    .c(al_944d9d4),
    .o({al_f373539a,al_c67bebad[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_edf2dc1f (
    .a(al_1315ed94[27]),
    .b(al_11033702[27]),
    .c(al_23e4bcdc),
    .o({al_45f4f2c6,al_c67bebad[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a98a3ed7 (
    .a(al_1315ed94[28]),
    .b(al_11033702[28]),
    .c(al_45f4f2c6),
    .o({al_ddde0c42,al_c67bebad[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_168d24d3 (
    .a(al_1315ed94[29]),
    .b(al_11033702[29]),
    .c(al_ddde0c42),
    .o({al_6fbb2d82,al_c67bebad[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c524c75b (
    .a(al_1315ed94[30]),
    .b(al_11033702[30]),
    .c(al_6fbb2d82),
    .o({al_a9d932ce,al_c67bebad[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86f90ba9 (
    .a(al_1315ed94[31]),
    .b(al_11033702[31]),
    .c(al_a9d932ce),
    .o({al_ecfcb3a4,al_c67bebad[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_344fb63e (
    .a(al_1315ed94[32]),
    .b(al_11033702[32]),
    .c(al_ecfcb3a4),
    .o({al_a3626bfc,al_c67bebad[32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fafc8f53 (
    .a(al_1315ed94[33]),
    .b(al_11033702[33]),
    .c(al_a3626bfc),
    .o({al_9031f908,al_c67bebad[33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33de60a (
    .a(al_1315ed94[34]),
    .b(al_11033702[34]),
    .c(al_9031f908),
    .o({al_94ad97ab,al_c67bebad[34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ae4de70 (
    .a(al_1315ed94[35]),
    .b(al_11033702[35]),
    .c(al_94ad97ab),
    .o({al_a6a5fe68,al_c67bebad[35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff46470e (
    .a(al_1315ed94[36]),
    .b(al_11033702[36]),
    .c(al_a6a5fe68),
    .o({al_467db6bc,al_c67bebad[36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68abff86 (
    .a(al_1315ed94[1]),
    .b(al_11033702[1]),
    .c(al_f373539a),
    .o({al_750066a4,al_c67bebad[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc96c084 (
    .a(al_1315ed94[37]),
    .b(al_11033702[37]),
    .c(al_467db6bc),
    .o({al_2c4eadf4,al_c67bebad[37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc93f476 (
    .a(al_1315ed94[38]),
    .b(al_11033702[38]),
    .c(al_2c4eadf4),
    .o({al_136010db,al_c67bebad[38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bea0d2b8 (
    .a(al_1315ed94[39]),
    .b(al_11033702[39]),
    .c(al_136010db),
    .o({al_3e351de0,al_c67bebad[39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_368990f0 (
    .a(al_1315ed94[40]),
    .b(al_11033702[40]),
    .c(al_3e351de0),
    .o({al_89cd14a1,al_c67bebad[40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ba912dab (
    .a(al_1315ed94[41]),
    .b(al_11033702[41]),
    .c(al_89cd14a1),
    .o({al_7e7ca026,al_c67bebad[41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a081c0b2 (
    .a(al_1315ed94[42]),
    .b(al_11033702[42]),
    .c(al_7e7ca026),
    .o({al_cde0b283,al_c67bebad[42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_458b8f4d (
    .a(al_1315ed94[43]),
    .b(al_11033702[43]),
    .c(al_cde0b283),
    .o({open_n3,al_c67bebad[43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_1315ed94[2]),
    .b(al_11033702[2]),
    .c(al_750066a4),
    .o({al_74601237,al_c67bebad[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_1315ed94[3]),
    .b(al_11033702[3]),
    .c(al_74601237),
    .o({al_9ea60d40,al_c67bebad[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_1315ed94[4]),
    .b(al_11033702[4]),
    .c(al_9ea60d40),
    .o({al_66e20fd7,al_c67bebad[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_1315ed94[5]),
    .b(al_11033702[5]),
    .c(al_66e20fd7),
    .o({al_c42610d7,al_c67bebad[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_1315ed94[6]),
    .b(al_11033702[6]),
    .c(al_c42610d7),
    .o({al_aafcdc4e,al_c67bebad[6]}));

endmodule 

