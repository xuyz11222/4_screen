// Verilog netlist created by Tang Dynasty v5.6.71036
// Sat Nov  2 12:33:56 2024

`timescale 1ns / 1ps
module div
  (
  clk,
  denominator,
  numerator,
  rst,
  start,
  done,
  quotient,
  remainder
  );

  input clk;
  input [11:0] denominator;
  input [26:0] numerator;
  input rst;
  input start;
  output done;
  output [26:0] quotient;
  output [11:0] remainder;

  parameter S_DEN = "UNSIGNED";
  parameter S_NUM = "UNSIGNED";
  parameter W_DEN = 12;
  parameter W_NUM = 27;
  // localparam W_CNT = 5;
  wire [4:0] al_1deac949;
  wire [4:0] al_d0dc52fd;
  wire [37:0] al_11033702;
  wire [37:0] al_1c1b24e7;
  wire [26:0] al_1315ed94;
  wire [26:0] al_9bfb1470;
  wire [37:0] al_c67bebad;
  wire [26:0] al_327525b3;
  wire al_a54c39e7;
  wire al_f74b2bbe;
  wire al_ea5880d3;
  wire al_bbe9aae2;
  wire al_d9ef6091;
  wire al_7109a3cd;
  wire al_f1bac0a6;
  wire al_61c118b2;
  wire al_9bb03b7;
  wire al_ea32c6e1;
  wire al_2ac97405;
  wire al_a0ebd25;
  wire al_f77a35ee;
  wire al_2902a00c;
  wire al_94925fa9;
  wire al_51a70210;
  wire al_fbeca432;
  wire al_ca5b12bc;
  wire al_b49c276a;
  wire al_a23af5a4;
  wire al_fe2986b6;
  wire al_875c79d9;
  wire al_d21ff3d4;
  wire al_20da7cd1;
  wire al_4b6c2990;
  wire al_2a9315a6;
  wire al_b9c5d958;
  wire al_56630a35;
  wire al_a1b0b17a;
  wire al_114eba31;
  wire al_c61b4192;
  wire al_d807637c;
  wire al_9993b324;
  wire al_1cfb05a7;
  wire al_6dd34b46;
  wire al_e5f94c1c;
  wire al_fec49048;
  wire al_610195b4;
  wire al_6d88e187;
  wire al_db08a961;
  wire al_9e273556;
  wire al_3e2f8c17;
  wire al_fc3d1d09;
  wire al_e7df159e;
  wire al_dd3ae65d;
  wire al_a2c118f2;
  wire al_738c830a;
  wire al_9ac6fc14;
  wire al_d35b5909;
  wire al_a6b4c38e;
  wire al_52a1be34;
  wire al_4edc63f3;
  wire al_1554169;
  wire al_f2c0d78d;
  wire al_52c3abfd;
  wire al_98a85355;
  wire al_d2d366b2;
  wire al_8ca46d3f;
  wire al_8fb8614f;
  wire al_bf599b52;

  AL_MAP_LUT6 #(
    .EQN("~(~A*~(~B*~(~C*(~(D)*~(E)*~(F)+D*E*F))))"),
    .INIT(64'hbabbbbbbbbbbbbba))
    al_f17cd423 (
    .a(start),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .e(al_1deac949[3]),
    .f(al_1deac949[4]),
    .o(al_d0dc52fd[0]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_147e6a1b (
    .a(start),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .o(al_d0dc52fd[1]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*~A)"),
    .INIT(32'h10000000))
    al_c8620855 (
    .a(al_1deac949[0]),
    .b(al_1deac949[1]),
    .c(al_1deac949[2]),
    .d(al_1deac949[3]),
    .e(al_1deac949[4]),
    .o(al_114eba31));
  AL_MAP_LUT5 #(
    .EQN("(~B*~A*(E@(D*C)))"),
    .INIT(32'h01111000))
    al_56322a5c (
    .a(al_114eba31),
    .b(start),
    .c(al_1deac949[0]),
    .d(al_1deac949[1]),
    .e(al_1deac949[2]),
    .o(al_d0dc52fd[2]));
  AL_MAP_LUT6 #(
    .EQN("(~A*(B*C*D*~(E)*~(F)+~(B)*~(C)*~(D)*E*~(F)+B*~(C)*~(D)*E*~(F)+~(B)*C*~(D)*E*~(F)+B*C*~(D)*E*~(F)+~(B)*~(C)*D*E*~(F)+B*~(C)*D*E*~(F)+~(B)*C*D*E*~(F)+B*C*D*~(E)*F+~(B)*~(C)*~(D)*E*F+B*~(C)*~(D)*E*F+~(B)*C*~(D)*E*F+B*C*~(D)*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F))"),
    .INIT(64'h1455400015554000))
    al_6614de08 (
    .a(start),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .e(al_1deac949[3]),
    .f(al_1deac949[4]),
    .o(al_d0dc52fd[3]));
  AL_MAP_LUT6 #(
    .EQN("(~A*(B*C*(E*D)*~(F)+~(B)*~(C)*~((E*D))*F+B*~(C)*~((E*D))*F+~(B)*C*~((E*D))*F+B*C*~((E*D))*F+B*~(C)*(E*D)*F+~(B)*C*(E*D)*F))"),
    .INIT(64'h1455555540000000))
    al_6dc5f615 (
    .a(start),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .e(al_1deac949[3]),
    .f(al_1deac949[4]),
    .o(al_d0dc52fd[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_cdf87825 (
    .a(denominator[0]),
    .b(start),
    .c(al_11033702[27]),
    .o(al_1c1b24e7[26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e6264f31 (
    .a(denominator[1]),
    .b(start),
    .c(al_11033702[28]),
    .o(al_1c1b24e7[27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_934b4c16 (
    .a(denominator[2]),
    .b(start),
    .c(al_11033702[29]),
    .o(al_1c1b24e7[28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_9fe68c39 (
    .a(denominator[3]),
    .b(start),
    .c(al_11033702[30]),
    .o(al_1c1b24e7[29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_41104578 (
    .a(denominator[4]),
    .b(start),
    .c(al_11033702[31]),
    .o(al_1c1b24e7[30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_12c43e12 (
    .a(denominator[5]),
    .b(start),
    .c(al_11033702[32]),
    .o(al_1c1b24e7[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_ded93226 (
    .a(denominator[6]),
    .b(start),
    .c(al_11033702[33]),
    .o(al_1c1b24e7[32]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_c35e0dcc (
    .a(denominator[7]),
    .b(start),
    .c(al_11033702[34]),
    .o(al_1c1b24e7[33]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_362a2d70 (
    .a(denominator[8]),
    .b(start),
    .c(al_11033702[35]),
    .o(al_1c1b24e7[34]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_619d59f3 (
    .a(denominator[9]),
    .b(start),
    .c(al_11033702[36]),
    .o(al_1c1b24e7[35]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8b9da26a (
    .a(denominator[10]),
    .b(start),
    .c(al_11033702[37]),
    .o(al_1c1b24e7[36]));
  AL_DFF_0 al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_114eba31),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_affc23c8 (
    .a(al_c61b4192),
    .b(numerator[0]),
    .c(start),
    .d(al_1315ed94[0]),
    .e(al_c67bebad[0]),
    .o(al_9bfb1470[0]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_7e4247d5 (
    .a(al_c61b4192),
    .b(numerator[10]),
    .c(start),
    .d(al_1315ed94[10]),
    .e(al_c67bebad[10]),
    .o(al_9bfb1470[10]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_8f76e334 (
    .a(al_c61b4192),
    .b(numerator[11]),
    .c(start),
    .d(al_1315ed94[11]),
    .e(al_c67bebad[11]),
    .o(al_9bfb1470[11]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_43c29c9e (
    .a(al_c61b4192),
    .b(numerator[12]),
    .c(start),
    .d(al_1315ed94[12]),
    .e(al_c67bebad[12]),
    .o(al_9bfb1470[12]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_dcb75b0 (
    .a(al_c61b4192),
    .b(numerator[13]),
    .c(start),
    .d(al_1315ed94[13]),
    .e(al_c67bebad[13]),
    .o(al_9bfb1470[13]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_e1773c9b (
    .a(al_c61b4192),
    .b(numerator[14]),
    .c(start),
    .d(al_1315ed94[14]),
    .e(al_c67bebad[14]),
    .o(al_9bfb1470[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_8e3693cb (
    .a(al_c61b4192),
    .b(numerator[15]),
    .c(start),
    .d(al_1315ed94[15]),
    .e(al_c67bebad[15]),
    .o(al_9bfb1470[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_79948be9 (
    .a(al_c61b4192),
    .b(numerator[16]),
    .c(start),
    .d(al_1315ed94[16]),
    .e(al_c67bebad[16]),
    .o(al_9bfb1470[16]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_cd0015f2 (
    .a(al_c61b4192),
    .b(numerator[17]),
    .c(start),
    .d(al_1315ed94[17]),
    .e(al_c67bebad[17]),
    .o(al_9bfb1470[17]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_5eba52cf (
    .a(al_c61b4192),
    .b(numerator[18]),
    .c(start),
    .d(al_1315ed94[18]),
    .e(al_c67bebad[18]),
    .o(al_9bfb1470[18]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_fd435063 (
    .a(al_c61b4192),
    .b(numerator[19]),
    .c(start),
    .d(al_1315ed94[19]),
    .e(al_c67bebad[19]),
    .o(al_9bfb1470[19]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_db832082 (
    .a(al_c61b4192),
    .b(numerator[1]),
    .c(start),
    .d(al_1315ed94[1]),
    .e(al_c67bebad[1]),
    .o(al_9bfb1470[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_e01dd5be (
    .a(al_c61b4192),
    .b(numerator[20]),
    .c(start),
    .d(al_1315ed94[20]),
    .e(al_c67bebad[20]),
    .o(al_9bfb1470[20]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_3caca9c9 (
    .a(al_c61b4192),
    .b(numerator[21]),
    .c(start),
    .d(al_1315ed94[21]),
    .e(al_c67bebad[21]),
    .o(al_9bfb1470[21]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_daadae89 (
    .a(al_c61b4192),
    .b(numerator[22]),
    .c(start),
    .d(al_1315ed94[22]),
    .e(al_c67bebad[22]),
    .o(al_9bfb1470[22]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_29e14add (
    .a(al_c61b4192),
    .b(numerator[23]),
    .c(start),
    .d(al_1315ed94[23]),
    .e(al_c67bebad[23]),
    .o(al_9bfb1470[23]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_144036ec (
    .a(al_c61b4192),
    .b(numerator[24]),
    .c(start),
    .d(al_1315ed94[24]),
    .e(al_c67bebad[24]),
    .o(al_9bfb1470[24]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_b86a6dbf (
    .a(al_11033702[12]),
    .b(al_11033702[13]),
    .c(al_11033702[14]),
    .d(al_1315ed94[12]),
    .e(al_1315ed94[13]),
    .f(al_1315ed94[14]),
    .o(al_d807637c));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(~C*A))"),
    .INIT(16'hc431))
    al_77e14fad (
    .a(al_11033702[23]),
    .b(al_11033702[24]),
    .c(al_1315ed94[23]),
    .d(al_1315ed94[24]),
    .o(al_fec49048));
  AL_MAP_LUT5 #(
    .EQN("(E*B*A*~(D@C))"),
    .INIT(32'h80080000))
    al_20244fba (
    .a(al_6dd34b46),
    .b(al_e5f94c1c),
    .c(al_11033702[22]),
    .d(al_1315ed94[22]),
    .e(al_fec49048),
    .o(al_610195b4));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    al_822ef4cd (
    .a(al_11033702[17]),
    .b(al_11033702[18]),
    .c(al_1315ed94[17]),
    .d(al_1315ed94[18]),
    .o(al_6d88e187));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    al_4609c472 (
    .a(al_6d88e187),
    .b(al_11033702[15]),
    .c(al_11033702[16]),
    .d(al_1315ed94[15]),
    .e(al_1315ed94[16]),
    .o(al_db08a961));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E)"),
    .INIT(32'h088cceef))
    al_bdafae35 (
    .a(al_11033702[13]),
    .b(al_11033702[14]),
    .c(al_1315ed94[12]),
    .d(al_1315ed94[13]),
    .e(al_1315ed94[14]),
    .o(al_9e273556));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((D*~A))*~(E)*~(F)+B*~(C)*~((D*~A))*~(E)*~(F)+~(B)*C*~((D*~A))*~(E)*~(F)+B*C*~((D*~A))*~(E)*~(F)+B*~(C)*(D*~A)*~(E)*~(F)+~(B)*C*(D*~A)*~(E)*~(F)+B*C*(D*~A)*~(E)*~(F)+B*~(C)*~((D*~A))*E*~(F)+~(B)*C*~((D*~A))*E*~(F)+B*C*~((D*~A))*E*~(F)+~(B)*C*(D*~A)*E*~(F)+B*C*(D*~A)*E*~(F)+~(B)*C*~((D*~A))*~(E)*F+B*C*~((D*~A))*~(E)*F+B*C*(D*~A)*~(E)*F+B*C*~((D*~A))*E*F)"),
    .INIT(64'h80c0e0f0f8fcfeff))
    al_7e9696d3 (
    .a(al_11033702[16]),
    .b(al_11033702[17]),
    .c(al_11033702[18]),
    .d(al_1315ed94[16]),
    .e(al_1315ed94[17]),
    .f(al_1315ed94[18]),
    .o(al_3e2f8c17));
  AL_MAP_LUT6 #(
    .EQN("(B*~(E*~A*~(C*~(F*D))))"),
    .INIT(64'h88c8ccccc8c8cccc))
    al_2f60b39a (
    .a(al_1cfb05a7),
    .b(al_610195b4),
    .c(al_db08a961),
    .d(al_9e273556),
    .e(al_3e2f8c17),
    .f(al_9993b324),
    .o(al_fc3d1d09));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_effa13b4 (
    .a(al_11033702[6]),
    .b(al_11033702[9]),
    .c(al_11033702[11]),
    .d(al_1315ed94[6]),
    .e(al_1315ed94[9]),
    .f(al_1315ed94[11]),
    .o(al_e7df159e));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_6dbdc742 (
    .a(al_11033702[8]),
    .b(al_11033702[10]),
    .c(al_1315ed94[8]),
    .d(al_1315ed94[10]),
    .o(al_dd3ae65d));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    al_e20893c3 (
    .a(al_e7df159e),
    .b(al_dd3ae65d),
    .c(al_11033702[7]),
    .d(al_1315ed94[7]),
    .o(al_a2c118f2));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_4be0c939 (
    .a(al_11033702[15]),
    .b(al_11033702[17]),
    .c(al_11033702[18]),
    .d(al_1315ed94[15]),
    .e(al_1315ed94[17]),
    .f(al_1315ed94[18]),
    .o(al_9993b324));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((~C*A))*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+~(B)*(~C*A)*D)"),
    .INIT(16'hf731))
    al_4718f307 (
    .a(al_11033702[0]),
    .b(al_11033702[1]),
    .c(al_1315ed94[0]),
    .d(al_1315ed94[1]),
    .o(al_f74b2bbe));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*C*D*E)"),
    .INIT(32'h40d0f4fd))
    al_c1df29b8 (
    .a(al_f74b2bbe),
    .b(al_11033702[2]),
    .c(al_11033702[3]),
    .d(al_1315ed94[2]),
    .e(al_1315ed94[3]),
    .o(al_738c830a));
  AL_MAP_LUT6 #(
    .EQN("(A*(~(B)*~(C)*~(D)*~(E)*~(F)+~(B)*~(C)*~(D)*E*~(F)+B*~(C)*~(D)*E*~(F)+~(B)*C*~(D)*E*~(F)+~(B)*~(C)*~(D)*~(E)*F+B*~(C)*~(D)*~(E)*F+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*~(C)*D*~(E)*F+~(B)*~(C)*~(D)*E*F+B*~(C)*~(D)*E*F+~(B)*C*~(D)*E*F+B*C*~(D)*E*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F))"),
    .INIT(64'h2aaa02aa002a0002))
    al_3e227b58 (
    .a(al_a2c118f2),
    .b(al_738c830a),
    .c(al_11033702[4]),
    .d(al_11033702[5]),
    .e(al_1315ed94[4]),
    .f(al_1315ed94[5]),
    .o(al_9ac6fc14));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((C*~A))*~(D)+B*~((C*~A))*~(D)+B*(C*~A)*~(D)+B*~((C*~A))*D)"),
    .INIT(16'h8cef))
    al_d3257d21 (
    .a(al_11033702[19]),
    .b(al_11033702[20]),
    .c(al_1315ed94[19]),
    .d(al_1315ed94[20]),
    .o(al_d35b5909));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6aae187d (
    .a(al_11033702[23]),
    .b(al_1315ed94[23]),
    .o(al_a6b4c38e));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*~(D)*~(E)*~(F)+~(A)*C*~(D)*~(E)*~(F)+A*C*~(D)*~(E)*~(F)+~(A)*~(C)*D*~(E)*~(F)+A*~(C)*D*~(E)*~(F)+~(A)*C*D*~(E)*~(F)+A*C*D*~(E)*~(F)+A*C*~(D)*E*~(F)+~(A)*~(C)*D*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*D*E*~(F)+A*~(C)*D*~(E)*F+~(A)*C*D*~(E)*F+A*C*D*~(E)*F+A*C*D*E*F))"),
    .INIT(64'h2000320033203332))
    al_12d215b6 (
    .a(al_d35b5909),
    .b(al_a6b4c38e),
    .c(al_11033702[21]),
    .d(al_11033702[22]),
    .e(al_1315ed94[21]),
    .f(al_1315ed94[22]),
    .o(al_52a1be34));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    al_cf5f85a (
    .a(al_11033702[24]),
    .b(al_11033702[25]),
    .c(al_1315ed94[24]),
    .d(al_1315ed94[25]),
    .o(al_4edc63f3));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_c1d3403 (
    .a(al_11033702[25]),
    .b(al_1315ed94[25]),
    .o(al_1554169));
  AL_MAP_LUT6 #(
    .EQN("(~((~D*~(C*~(B*~A))))*~(E)*~(F)+~((~D*~(C*~(B*~A))))*E*~(F)+(~D*~(C*~(B*~A)))*E*~(F)+~((~D*~(C*~(B*~A))))*E*F)"),
    .INIT(64'hffb00000ffffffb0))
    al_967c6e26 (
    .a(al_52a1be34),
    .b(al_fec49048),
    .c(al_4edc63f3),
    .d(al_1554169),
    .e(al_11033702[26]),
    .f(al_1315ed94[26]),
    .o(al_f2c0d78d));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_be651df4 (
    .a(al_11033702[6]),
    .b(al_1315ed94[6]),
    .o(al_a54c39e7));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6db3ef19 (
    .a(al_11033702[9]),
    .b(al_1315ed94[9]),
    .o(al_52c3abfd));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    al_115bf27e (
    .a(al_d807637c),
    .b(al_9993b324),
    .c(al_11033702[16]),
    .d(al_1315ed94[16]),
    .o(al_1cfb05a7));
  AL_MAP_LUT6 #(
    .EQN("(~B*(~(A)*~(C)*~(D)*~(E)*~(F)+~(A)*C*~(D)*~(E)*~(F)+A*C*~(D)*~(E)*~(F)+~(A)*~(C)*D*~(E)*~(F)+A*~(C)*D*~(E)*~(F)+~(A)*C*D*~(E)*~(F)+A*C*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+~(A)*~(C)*D*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*D*E*~(F)+~(A)*~(C)*D*~(E)*F+~(A)*C*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*D*E*F))"),
    .INIT(64'h1000310033103331))
    al_d40072f7 (
    .a(al_a54c39e7),
    .b(al_52c3abfd),
    .c(al_11033702[7]),
    .d(al_11033702[8]),
    .e(al_1315ed94[7]),
    .f(al_1315ed94[8]),
    .o(al_98a85355));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9b8487df (
    .a(al_11033702[9]),
    .b(al_1315ed94[9]),
    .o(al_d2d366b2));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+~((~B*~A))*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+(~B*~A)*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*C*D*E*F)"),
    .INIT(64'he000fe00ffe0fffe))
    al_75242fbe (
    .a(al_98a85355),
    .b(al_d2d366b2),
    .c(al_11033702[10]),
    .d(al_11033702[11]),
    .e(al_1315ed94[10]),
    .f(al_1315ed94[11]),
    .o(al_8ca46d3f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_2f9da10c (
    .a(al_11033702[31]),
    .b(al_11033702[32]),
    .c(al_11033702[33]),
    .d(al_11033702[34]),
    .e(al_11033702[35]),
    .f(al_11033702[36]),
    .o(al_8fb8614f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_90c42bd9 (
    .a(al_8fb8614f),
    .b(al_11033702[27]),
    .c(al_11033702[28]),
    .d(al_11033702[29]),
    .e(al_11033702[30]),
    .f(al_11033702[37]),
    .o(al_bf599b52));
  AL_MAP_LUT6 #(
    .EQN("(F*~(C*~(A*~(E*D*~B))))"),
    .INIT(64'h8fafafaf00000000))
    al_6b244534 (
    .a(al_fc3d1d09),
    .b(al_9ac6fc14),
    .c(al_f2c0d78d),
    .d(al_8ca46d3f),
    .e(al_1cfb05a7),
    .f(al_bf599b52),
    .o(al_c61b4192));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_f30062e5 (
    .a(al_c61b4192),
    .b(numerator[25]),
    .c(start),
    .d(al_1315ed94[25]),
    .e(al_c67bebad[25]),
    .o(al_9bfb1470[25]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_7378e3a9 (
    .a(al_11033702[19]),
    .b(al_11033702[20]),
    .c(al_11033702[21]),
    .d(al_1315ed94[19]),
    .e(al_1315ed94[20]),
    .f(al_1315ed94[21]),
    .o(al_6dd34b46));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_6c1e3994 (
    .a(al_11033702[25]),
    .b(al_11033702[26]),
    .c(al_1315ed94[25]),
    .d(al_1315ed94[26]),
    .o(al_e5f94c1c));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_47ac1c09 (
    .a(al_c61b4192),
    .b(numerator[26]),
    .c(start),
    .d(al_1315ed94[26]),
    .e(al_c67bebad[26]),
    .o(al_9bfb1470[26]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_3e04c0e7 (
    .a(al_c61b4192),
    .b(numerator[2]),
    .c(start),
    .d(al_1315ed94[2]),
    .e(al_c67bebad[2]),
    .o(al_9bfb1470[2]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_b86e3fac (
    .a(al_c61b4192),
    .b(numerator[3]),
    .c(start),
    .d(al_1315ed94[3]),
    .e(al_c67bebad[3]),
    .o(al_9bfb1470[3]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_1f499def (
    .a(al_c61b4192),
    .b(numerator[4]),
    .c(start),
    .d(al_1315ed94[4]),
    .e(al_c67bebad[4]),
    .o(al_9bfb1470[4]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_8f1711f3 (
    .a(al_c61b4192),
    .b(numerator[5]),
    .c(start),
    .d(al_1315ed94[5]),
    .e(al_c67bebad[5]),
    .o(al_9bfb1470[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_6e1c653d (
    .a(al_c61b4192),
    .b(numerator[6]),
    .c(start),
    .d(al_1315ed94[6]),
    .e(al_c67bebad[6]),
    .o(al_9bfb1470[6]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_b46e3fd7 (
    .a(al_c61b4192),
    .b(numerator[7]),
    .c(start),
    .d(al_1315ed94[7]),
    .e(al_c67bebad[7]),
    .o(al_9bfb1470[7]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_d21f8608 (
    .a(al_c61b4192),
    .b(numerator[8]),
    .c(start),
    .d(al_1315ed94[8]),
    .e(al_c67bebad[8]),
    .o(al_9bfb1470[8]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*B*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B*C)"),
    .INIT(32'hcfcac5c0))
    al_42e41119 (
    .a(al_c61b4192),
    .b(numerator[9]),
    .c(start),
    .d(al_1315ed94[9]),
    .e(al_c67bebad[9]),
    .o(al_9bfb1470[9]));
  AL_DFF_0 al_b26d62bf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[0]));
  AL_DFF_0 al_809f7104 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[1]));
  AL_DFF_0 al_c1468025 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[2]));
  AL_DFF_0 al_c19d8344 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[3]));
  AL_DFF_0 al_ca1eda73 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[4]));
  AL_DFF_0 al_b40e8e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[8]));
  AL_DFF_0 al_2259e8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[9]));
  AL_DFF_0 al_5f624aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[10]));
  AL_DFF_0 al_d532b054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[11]));
  AL_DFF_0 al_9d987fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[12]));
  AL_DFF_0 al_220744cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[13]));
  AL_DFF_0 al_e241f44a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[14]));
  AL_DFF_0 al_897da5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[15]));
  AL_DFF_0 al_9e863954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[16]));
  AL_DFF_0 al_a186fcad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[17]));
  AL_DFF_0 al_fd544ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[0]));
  AL_DFF_0 al_21ba363c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[18]));
  AL_DFF_0 al_c602bc36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[19]));
  AL_DFF_0 al_be443a52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[21]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[20]));
  AL_DFF_0 al_961a8bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[22]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[21]));
  AL_DFF_0 al_6d594c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[23]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[22]));
  AL_DFF_0 al_5e95843a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[24]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[23]));
  AL_DFF_0 al_d701a9b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[25]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[24]));
  AL_DFF_0 al_420d26fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[26]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[25]));
  AL_DFF_0 al_eb274ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[26]));
  AL_DFF_0 al_59566ddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[27]));
  AL_DFF_0 al_40ebe0d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[1]));
  AL_DFF_0 al_88ac72e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[28]));
  AL_DFF_0 al_415d213a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[29]));
  AL_DFF_0 al_2589b38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[30]));
  AL_DFF_0 al_d3625316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[31]));
  AL_DFF_0 al_a773e9fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[32]));
  AL_DFF_0 al_b5a98930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[33]));
  AL_DFF_0 al_84e187a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[34]));
  AL_DFF_0 al_f3095820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[35]));
  AL_DFF_0 al_9b82a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[36]));
  AL_DFF_0 al_e2ab1094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[11]),
    .en(1'b1),
    .sr(~start),
    .ss(1'b0),
    .q(al_11033702[37]));
  AL_DFF_0 al_b4cd3408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[2]));
  AL_DFF_0 al_16607eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[3]));
  AL_DFF_0 al_2e1082f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[4]));
  AL_DFF_0 al_806f02ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[5]));
  AL_DFF_0 al_e97bb64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[6]));
  AL_DFF_0 al_f7f2da08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[7]));
  AL_DFF_0 al_596b0fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[8]));
  AL_DFF_0 al_5cfa2c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[9]));
  AL_DFF_0 al_c56c02f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[10]));
  AL_DFF_0 al_60ec2662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[11]));
  AL_DFF_0 al_ea3f598e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[12]));
  AL_DFF_0 al_dd4ae85d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[13]));
  AL_DFF_0 al_e2aa8055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[14]));
  AL_DFF_0 al_82aa8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[15]));
  AL_DFF_0 al_7f911c70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[16]));
  AL_DFF_0 al_8908ba38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[17]));
  AL_DFF_0 al_16ad90bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[0]));
  AL_DFF_0 al_2149b062 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[18]));
  AL_DFF_0 al_56d82898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[19]));
  AL_DFF_0 al_c8bec57f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[20]));
  AL_DFF_0 al_1f071837 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[21]));
  AL_DFF_0 al_9acbb644 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[22]));
  AL_DFF_0 al_286bd0de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[23]));
  AL_DFF_0 al_7e8bb9f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[24]));
  AL_DFF_0 al_d4e324dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[25]));
  AL_DFF_0 al_bcaf406d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[26]));
  AL_DFF_0 al_e1044ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[1]));
  AL_DFF_0 al_16da6de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[2]));
  AL_DFF_0 al_e819e904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[3]));
  AL_DFF_0 al_4990808d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[4]));
  AL_DFF_0 al_d51e17ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[5]));
  AL_DFF_0 al_b67f884b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[6]));
  AL_DFF_0 al_ff3308ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[7]));
  AL_DFF_0 al_c1e3ea45 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[8]));
  AL_DFF_0 al_b7aa029f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[9]));
  AL_DFF_0 al_2f4f18cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[10]));
  AL_DFF_0 al_42a7eb97 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[11]));
  AL_DFF_0 al_f77c099a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[12]));
  AL_DFF_0 al_6893ba8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[13]));
  AL_DFF_0 al_d6d1e991 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[14]));
  AL_DFF_0 al_4d3bf6cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[15]));
  AL_DFF_0 al_aa8c310 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[16]));
  AL_DFF_0 al_d8095998 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[17]));
  AL_DFF_0 al_53efe64b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[0]));
  AL_DFF_0 al_68082bd4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[18]));
  AL_DFF_0 al_d9e8ef9f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[19]));
  AL_DFF_0 al_39169fb8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[20]));
  AL_DFF_0 al_c179532 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[21]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[21]));
  AL_DFF_0 al_7d105784 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[22]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[22]));
  AL_DFF_0 al_573a0a58 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[23]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[23]));
  AL_DFF_0 al_d0deffcb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[24]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[24]));
  AL_DFF_0 al_150254f9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[25]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[25]));
  AL_DFF_0 al_47f1ba67 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[26]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[26]));
  AL_DFF_0 al_26890f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[1]));
  AL_DFF_0 al_802c7023 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[2]));
  AL_DFF_0 al_9c45670 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[3]));
  AL_DFF_0 al_b0a0e999 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[4]));
  AL_DFF_0 al_739d9f2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[5]));
  AL_DFF_0 al_7f9eee7d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[6]));
  AL_DFF_0 al_741313a7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[7]));
  AL_DFF_0 al_ce6e5997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[8]));
  AL_DFF_0 al_7c322425 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[9]));
  AL_DFF_0 al_1f65ec13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[10]));
  AL_DFF_0 al_63457b5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[11]));
  AL_DFF_0 al_11fe6cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[12]));
  AL_DFF_0 al_9cfb6f54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[13]));
  AL_DFF_0 al_40b705d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[14]));
  AL_DFF_0 al_cbb21b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[15]));
  AL_DFF_0 al_a743530c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[16]));
  AL_DFF_0 al_50032887 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[17]));
  AL_DFF_0 al_5e904a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c61b4192),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[0]));
  AL_DFF_0 al_db3b2b53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[18]));
  AL_DFF_0 al_4496adb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[19]));
  AL_DFF_0 al_db38e2c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[20]));
  AL_DFF_0 al_b910420c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[21]));
  AL_DFF_0 al_90d7e42b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[21]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[22]));
  AL_DFF_0 al_f16a60a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[22]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[23]));
  AL_DFF_0 al_91adf23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[23]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[24]));
  AL_DFF_0 al_77ecd5d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[24]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[25]));
  AL_DFF_0 al_149f3658 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[25]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[26]));
  AL_DFF_0 al_116f1db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[1]));
  AL_DFF_0 al_6c993e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[2]));
  AL_DFF_0 al_23963ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[3]));
  AL_DFF_0 al_6c25cf29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[4]));
  AL_DFF_0 al_e7cc423c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[5]));
  AL_DFF_0 al_2c6ea385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[6]));
  AL_DFF_0 al_a356779f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[7]));
  AL_DFF_0 al_f27b108d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[8]));
  AL_DFF_0 al_d1a67c2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[9]));
  AL_DFF_0 al_a7f95d18 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[10]));
  AL_DFF_0 al_da9c9cea (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[11]));
  AL_DFF_0 al_cbbb4490 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[0]));
  AL_DFF_0 al_30153836 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[1]));
  AL_DFF_0 al_37ead40d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[2]));
  AL_DFF_0 al_7625712c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[3]));
  AL_DFF_0 al_2531de5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[4]));
  AL_DFF_0 al_2ccbdc6d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[5]));
  AL_DFF_0 al_2c62c395 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[6]));
  AL_DFF_0 al_ee1990ef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_1315ed94[7]),
    .b(al_11033702[7]),
    .c(al_ea32c6e1),
    .o({al_2ac97405,al_c67bebad[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_1315ed94[8]),
    .b(al_11033702[8]),
    .c(al_2ac97405),
    .o({al_a0ebd25,al_c67bebad[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_1315ed94[9]),
    .b(al_11033702[9]),
    .c(al_a0ebd25),
    .o({al_f77a35ee,al_c67bebad[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_1315ed94[10]),
    .b(al_11033702[10]),
    .c(al_f77a35ee),
    .o({al_2902a00c,al_c67bebad[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_1315ed94[11]),
    .b(al_11033702[11]),
    .c(al_2902a00c),
    .o({al_94925fa9,al_c67bebad[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_1315ed94[12]),
    .b(al_11033702[12]),
    .c(al_94925fa9),
    .o({al_51a70210,al_c67bebad[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_1315ed94[13]),
    .b(al_11033702[13]),
    .c(al_51a70210),
    .o({al_fbeca432,al_c67bebad[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_1315ed94[14]),
    .b(al_11033702[14]),
    .c(al_fbeca432),
    .o({al_ca5b12bc,al_c67bebad[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_1315ed94[15]),
    .b(al_11033702[15]),
    .c(al_ca5b12bc),
    .o({al_b49c276a,al_c67bebad[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_1315ed94[16]),
    .b(al_11033702[16]),
    .c(al_b49c276a),
    .o({al_a23af5a4,al_c67bebad[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f5224f5b (
    .a(1'b0),
    .o({al_ea5880d3,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_1315ed94[17]),
    .b(al_11033702[17]),
    .c(al_a23af5a4),
    .o({al_fe2986b6,al_c67bebad[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bbcbdbe (
    .a(al_1315ed94[18]),
    .b(al_11033702[18]),
    .c(al_fe2986b6),
    .o({al_875c79d9,al_c67bebad[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_216ec453 (
    .a(al_1315ed94[19]),
    .b(al_11033702[19]),
    .c(al_875c79d9),
    .o({al_d21ff3d4,al_c67bebad[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c943a4d2 (
    .a(al_1315ed94[20]),
    .b(al_11033702[20]),
    .c(al_d21ff3d4),
    .o({al_20da7cd1,al_c67bebad[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_920ee641 (
    .a(al_1315ed94[21]),
    .b(al_11033702[21]),
    .c(al_20da7cd1),
    .o({al_4b6c2990,al_c67bebad[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e359bb16 (
    .a(al_1315ed94[22]),
    .b(al_11033702[22]),
    .c(al_4b6c2990),
    .o({al_2a9315a6,al_c67bebad[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a6af83b3 (
    .a(al_1315ed94[23]),
    .b(al_11033702[23]),
    .c(al_2a9315a6),
    .o({al_b9c5d958,al_c67bebad[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_717da7cc (
    .a(al_1315ed94[24]),
    .b(al_11033702[24]),
    .c(al_b9c5d958),
    .o({al_56630a35,al_c67bebad[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_916a9569 (
    .a(al_1315ed94[25]),
    .b(al_11033702[25]),
    .c(al_56630a35),
    .o({al_a1b0b17a,al_c67bebad[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b53f57fa (
    .a(al_1315ed94[26]),
    .b(al_11033702[26]),
    .c(al_a1b0b17a),
    .o({open_n3,al_c67bebad[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6e3dfcf (
    .a(al_1315ed94[0]),
    .b(al_11033702[0]),
    .c(al_ea5880d3),
    .o({al_bbe9aae2,al_c67bebad[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68abff86 (
    .a(al_1315ed94[1]),
    .b(al_11033702[1]),
    .c(al_bbe9aae2),
    .o({al_d9ef6091,al_c67bebad[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_1315ed94[2]),
    .b(al_11033702[2]),
    .c(al_d9ef6091),
    .o({al_7109a3cd,al_c67bebad[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_1315ed94[3]),
    .b(al_11033702[3]),
    .c(al_7109a3cd),
    .o({al_f1bac0a6,al_c67bebad[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_1315ed94[4]),
    .b(al_11033702[4]),
    .c(al_f1bac0a6),
    .o({al_61c118b2,al_c67bebad[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_1315ed94[5]),
    .b(al_11033702[5]),
    .c(al_61c118b2),
    .o({al_9bb03b7,al_c67bebad[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_1315ed94[6]),
    .b(al_11033702[6]),
    .c(al_9bb03b7),
    .o({al_ea32c6e1,al_c67bebad[6]}));

endmodule 

