

module hdmi_tx_controller_wrapper #(
    parameter HTOTAL  = 2200,
    parameter HSA     = 44,
    parameter HFP     = 88,
    parameter HBP     = 148,
    parameter HACTIVE = 1920,
    parameter VTOTAL  = 1125,
    parameter VSA     = 5,
    parameter VFP     = 4,
    parameter VBP     = 36,
    parameter VACTIVE = 1080,

    parameter VIDEO_TPG = "Enable",

    parameter VIDEO_FORMAT      = "RGB444",
    parameter VIDEO_VIC         = 16,
    parameter AUDIO_CTS         = 148500,
    parameter AUDIO_N           = 6144,
    parameter AUDIO_SAMPLE_RATE = "48K"
)    
(
    input wire       I_pixel_clk,
    input wire       I_rst,

///**********************  video stream input  ***************************
    input wire       I_video_in_user,
    input wire       I_video_in_valid,
    input wire       I_video_in_last,
    input wire[23:0] I_video_in_data,
    output wire      O_video_in_ready,

///*********************  audio stream input  ***************************
    input wire       I_audio_valid,     
    input wire[23:0] I_audio_left_data, 
    input wire[23:0] I_audio_right_data,

///*********************  tmds data output  *****************************
    output wire[9:0] O_ch0_tmds_code_data,     
    output wire[9:0] O_ch1_tmds_code_data,     
    output wire[9:0] O_ch2_tmds_code_data,     
    output wire[9:0] O_clk_tmds_code_data      

);


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
k7Vs2r+Kqq6ituoNGbcbFi86smdG+Wibg94qT3NIumVw5lhBjDRM9FNmq9Zlonuy
PWWI4JdUsqCCtCJ0LgnbX0/xOHdwEPTy50dHdd1FCcdvmyyV1oND8p1zBz30SN7E
We609maEoS6APuD1e6oFveR/DTzLjXeUp2jrDhUyzuc=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 108528)
`pragma protect data_block
a1NGakdObHhFT1hkZFpXd6Jv3z4mv4k/6+tD2x+wR1QIX9vvnxnEZeOwZ8TwZcYJ
Rh2R1gaJ+l1jYnOdepnuzbZzVP1f8gGP6p15cSy6yFP6V8NcgWS+SVDI/HK/IvGh
oJ8eo2XjtbDOQBuPmSQ5QvhGv79BEChJqyCCcKqEIhNXKXvSaWYWSF/8w2aMYr8g
wvBpUhSr4H3zIEO9JH3g3v/q2oWAHZww29gKni3uBtq17r1Aj4UXKl+PZAbkQQ5W
4wuu2+ElyEfV4R7FxSxEiupJurdlZ8nKxfMu4V3MgY3iW3T6MNec8tOSluX6I4Rw
oORCAHwwEDZhtkJy4s7UeATBzTrRXqumr8qfAi27lZV2s0pGIbYHkBTkUWc6JXiY
nvEDgElFjNfksVqEj68VTD89480yo/lwUOmqglD1s5/h2SFOr1R31obMoy7JPTfZ
YSpC8Qrp9Tab8oIlEoyFeaaHARAr8Xvnn6+EA6PS9WxoYfB1LmFR/sWEZ8Jms/rq
RCP+1GYU5VmIZBZb9SjH09UOHjf+NfmX1s5HO7Qg4SMLCsyb3ZdRaamjhqWcDC3R
i6+ypsSRK8vdJpZwt8JA65ZM6+J6WTZmCud5FG6hoxmIl8WDW1QNDc2Ze/rhvnjc
4qDKSBBZowxTw3olcVqS9jQD9iLCgPrGerhyAEfXdWNliVfBzbpswVsWhK2cW2B1
Ozx807MilRs3oLSAayIaDOKkXTPTiLzu9aKStpph+ABiuzaVgrwU38hup6B1hjWL
SzWXt+eMqOyc7bAqyVDXI6tPYTp8zyiekNT3sP+bbIuUdpvXMw52dE6zLJFZK24d
yF/O6SjPvr6DeIChLDhb392RIdS5PBp1M40kwtIhgn1QUzNzJBPYkl+neHyXy+ib
uANbv24pT7GKBkS+Gu3ReHQZjmi0HLl4BWCx6AspYKUYH8G84L93UbEbKiZrdNRz
QgiRMQ0D5lWmYhtm03VAuQapY+fp5n07R5xdUUMSHJSxNftBw9QD6geR0cOTrQoZ
M4dEBMWyn2kh+ChY6ZlFQ6r9838D36H+iPIMjv/8XV4vQG5CvnzTTzfM9sueRVFW
CwdZK84L/0xPPhcrSsEYCD/GmT1n5JUCJ6wryXvwmOYk1U9eRGK0/gSHFIN8+7o+
bpYqiFMJYKoJ84PGYTdnX40FBLkIWOnVhst8BbR9UycNKnQh2xiFq3Q1xYMhUww7
zpnFkssPWIc5Ndnf7zckvVUx0TxzH7V9KjInpkqJ8fgbbsxaCDEuM1MnNLvJmV1W
XNpbq+eo1DlBgogBmvfCqnm4p/lNfC9IGEG9hK/GOb4G2SJrI7PZ2PZUHHh34bln
00eTHK1zDG7mCfeuCr/tjYHouzbzWjZSCma/8ckif8pn6wgZDTwzRSrgm4wOdjJK
f7A0KjdMg3NBz/kn3KkuCaTvWhQsLN73W9v0zJd1A8fkLvJbWH6D5njEmWteoQzW
LrKjIxarNVAr/3vNRfz6RxC+2Him3XBqUjmfzjyPTRsaAHc2oZRM50BB8Y/Itubi
GsNHYDTzfAZA+F2y4Tezfo9wTeg1Yu1PQYabMgbEgPQ0zPsqD9TW4BIqhlC44EAN
8eYxQrcJKBntONguNKxMS8wZyGClwFdRG9OPhmWsDNyUq6gMLHnAtYQEwisnTxAv
Eny6YltIZ/7UfzlQPln10/iT7qXQ3ld2T/1Gkih/qH2dl/pCno1xPPrYmOufXao5
PUzAwkYPCkVgzH4ojSVsSvTW3ShZigAQg3KmJ8ioqZ9yulvAhik/EWj1KkPUXWJI
kwlp1V+/jKvLAqJbCnfYbZHrFlR3MHycs4YzTQLUBVaxs8Sd3AQd5XMEOk8bsrcH
Cgl1AfXHqUX0oNEFChlH+hd6UHiE1/39BBpcEPjf9tolfLTUmY0cXCXTx/uxR+Tm
d8Q1sBMwiXN8fsE0xr454eIo3ov5//3OGDSP3TbsjnY6O0bIsuf58iNGFNUal7NC
NKSXALnS4H2sO4hhOCYp4BUmrjT1TTeDkSAE/Or0AOqLF4HQ7zR13EDMTshbxGll
DUk9ZKHsmxOgKmGFOL18MuP2wwgU/bEB2i30gct1prEv6lWphbJ5Vd8QivfLW9MF
yIfHJUzISwCRd7XzJhP8iIplzqNwdKRXWcHyD3e6+ErwNDQHrQVI7fMLJpRnuah3
XE+yeaOKVcwqu/Eyg3PMZvJyPDx3XlNpwxT92zm/wuKlFbMbCU+s/j6Q/layODx4
P4uv5ygbzbffX9B6JDHZ/Jj0NaPtH1voIqVh9HfGxAzLnU7mItQFLDeQM2iy4URI
TMRDuW4ptyxyVEOzQ2kFVxfFQ3hwGl7isigGCBqfn8/judlKLr0T/TOyA3IW8D4e
Lzpg0UBoVUZ40AeA4tdhRdNTRrmQHNa1udVD6t1cBP8JhqOaDeOGv+wc66X4+lVG
baX8xHsEA3E5R7OqSxMmIZT29we+sn3PW7QHkoVYefBgXgkQM/58r27gNiJRKENt
T5J/Y6RFJSC5yw96NKQpk0maXAPFRZv9BNkfTnEow5Is9pu+paya37QGulQQ4tdR
29vInCvVUBvpqwNpdqmKKSPdVvb1DCuKMlQMoqpWATKTM0XQoDlp8Y0nI81TdHWX
JPAhJhiQJ7xfyaCGHZyZW7rZ3Mq1CXxMZURzrDI4A7Ym4HJvakaJTIITcyzduk/k
r44uI7tM597UEikEaUF89s3PzbBmx3BOxM8rhQByvsctHHGuELux0jgLTogthmNT
xF2PZRL9E2jnXg0HkKTqRLTzYppF/wUVqiNVZs8qniWf7px2SEjOqPNYNubDqIM8
B1ItUL+kQkxc9VZUoqaGxZJFp5O9eqXuiWHolovwSvkp9ZbdYjDg8S+9TgltSVZn
LjPG1Y5lkannYYtuUjSWmwRjnyp6efaxXEIifo5+8Ka9lTqsoe0Z4xn61qYwQcIv
LqlS4KJT7Zaf4nu4AzhSbl4I7Wi7aicqSTXInCEyDATW+POguDjuwMBOILyFghxQ
ZxIcP/TwKzDi0/+a/zJDV5WTC5IaHNAU5Objgoe6Ik78jMtE6YIZI2pmFhfQ8LEb
dPfFutb7bOUTcJReAMPXebPZm9b35lY9bjfwUs391SxYKoyhwipQId1WPL1k2DYJ
XP6ASrWWwaEI1UhmVW3bXu54x+moJviWv3DDAbPvGoUPjKZJUoJTOE50BQWMbOnE
bJsbpNam2GjXDG7CNc0uiMoB9SVD2AYIEqf00DP4JUO2Lsh6W/6SowDusIfAZrHM
xsFQFsnp4L1P9qxjcGfxvcHLz11ezDzJGyOsZH7WVQ4x9Nzdkr2b5RqDmR4pG3Hz
8PMWqUuoArcTP4YujV9uzewLGxPdNcFOjpEgOrUs5ONRWEsBxB+D15ZBrZ/wSQq7
/9CkBDNDJ4fUyTNAdGfXOYg6m05att4Bi4bGHFR7q/FDq+xVbUjNrdxIW5uK/2hJ
WQKsNeWGzLLIAdl72H8KiCeQy3bbdJpRpQhtrcnJ5BtFF2cMCTZ7ayaYqav8Dnyp
oG7OKWLutcpSjTcl9ivn88DRjLHcmjc2B4ZfROj4ccXXEgJrveUF/aIVwpw7hJYR
RcWL6R6zY7KJbKreLyQeDMJ9kOF1dIVwRxM2doQ+DrtMLlsfjC+q/w+Ke/G8wwrf
PEchRD97RGOFuKYu7Tgb99lSEU6lr3R0pdKE5UVNV/o4PFNLC/zScOFzyE+CAQpV
oRJs+QiBcrk8IG13UpxPjuqfXHkqtbgAAU/RsYkh4Ql5YFd2wglCS73chnKiEU05
c8wb+utdOctZgNu9e15oMZ3oL/Bg58Ab2wXyi6oPRKkKvNzT4YLYgj/KlAbykowX
cVQJJUSNqob34iw3+4dhnf9vZpbZJGtqpANdL2I+/QzVTGumBxqydtXSdP9JU3ty
ja6LT0I/iO8iLEwUdyuReSB1xM00fGQhTDIgv+IItDHv+tgPI5IlR/cVOCizDApX
IZCsc5N8MK9iy4rSY9g0hMJeNRIfTEZdwqV3bP7Ex0SxpzIQINd7UGa37sV/1pEv
5cdIW75k4frLYdevgnYNi2uOazNQv1/nRjmiJOAFT1YBGx/IbkSzm+UuA9W2/jsH
WxYgLQo2oavletKA2U2VBIo5GP/jC5iIDmOQxMlgd/0P/U3CMHg5L1nVd93eEobt
sdLXX/P1vWKTki997oP9fuIR2KzettBOxo9pLVBcYyUkERTW0WTQVoBFnhH+Y/iZ
6w7rViplBShQ4zfPWGdths7GKofWW99JvUItBJDbL1ztqL6S3rQI3yMdOggrGzDj
SVTkFqSm7XZkF+JAmKOiuWKcWyMZ6awVZ1fi7gDSSi4Er7WsW4aY2rLzhAZmvfVB
IuaY9pVJay3WzyREjRGVfutxYSbhC6+W5TWOW8gqOFTyA8i8GY0S7ogjvz/XEuxq
/KbENs33dvbVk0+/ZhHn613jte0g1vNa5YoQjwqph2lC5v98Txw+Yx7wXSmSsX1H
SPy/rSWnsMVnwevwnJugE9aNOIvZq71Lc5gVoxEXCOOaIgFUixJidI1f6+O46NTW
JTuUP+mostl52vNQY6IWV6Dxef+UsFCwx2vY983RK4lO8X8UlunBX8LZp7qc4qiM
SVa0ogzVT/kMadMKZgrG5Uyw77jeo69E78ROgoxT2SBQvv+b2VBiW7jHHvemLQYd
m7D5QDqPZYXk2BFL22O1oIH3xuG+er0g1R//Xy0Zr1Ld2v1Kh1KldYF6MFrsLkyx
pcSupn13BtkV32VsaHckj6PH/oD0qXKHDGFiagaofuSAk8Wz9FHOAMdK/Zn0MFaR
EiO1ijcFUoZGdc8h1uui+6A3NydPHNinUtCV3v/E2u2HKK/WFMZ8PlajDhT097Xl
Vp/nls9ps0TWq1KZjaXpPG71rgmcMtOn1HbTNiTSQ3rkxli/x1m7hK22WrBNostj
2AgqirgoCbWVxbHektrwxw4svulbmymDWq6iE39y9IvJN0JGtNZH9CGR06xxe+bU
KIZYaQlkLxzHqc6mNQpL/cmIfPmArTKicyeh+mipLjp2HRXlxEaYZDi7pGEYkFyh
FlTyXH5sLEtm3XjxLi57NKXq9KQtI8hF0DoD8aQ1oCHihlSRfLT5xF7NSDu16Z1n
WWXh6Y9s5VjvRxZzR5zJ6FBAyRWOrO/7XYxxPNVRQnnaHxC6cB6vagWX+qit5kcj
ckIpcWSbgEuyPAzetAsznypsKf4L+Liqymb9KxSwkF1xajDP8NSugMRNPpc4+hEF
yIj0k9XOB3O9cqOlro/E1oCQjQJTkoCUtIGUC2kF4tCi/vjFCqdjIUnKgoJShG1G
D0GMV0xO5hYOwMcpH3/uFHIi349nTftrqDmFiMzWMF8sWfxxLD8KJnNuefJ9brHQ
ucsVmIEfV9wOcCvx155R8X+MmKCZjg+NXzzQXp+Xj/cpNuHQUywThBUvEIdviq2y
83Gn3C3t2dfLbjZnnym5Lyfi6aoL8SFbh6XJ3iwcQmkz8jzkkupqNEcf33+jS1uv
4MHgipn/lMGUQwHyrRMzt14CY5o8jMxESLFYf6cxG6C0bwifP3HdEMutaAuAp5lz
2WKpGKW88ziR6SIXOr0F/JbAHCBAbYXAFoq4QhfjAWJGZqbRXqZv1rZLFPvZUcxl
thqjZEDBrr06Fbyfa87edF9BoQV5K9CtN9RLgniohqZ6f7zBcaIly7OyZaIzywIC
3wfkiOOhB7URxUjtjaWpOV6+PzY10v3knmRjYgJp2L5vC1MfZOei2cZS7GRD2tug
KHKiZJx/lL84Uy7vlxxQZpUQ+Wmy/DMxH5L+IBKe+6tn1wlghtjbxNSDgoDy1iJy
LnBCE/Vu1L83DmKI39kw1iinzzk7Vk/r7SvB7Cc8INJ5dDbQZ7U3xH3/n503jy5R
rXTkxWEx6dIx8d7CfknKRWH74timnLCMT3b6IEft3WBLrS+Bdz6SwqeiPcbMms0Z
N1Vzdm2t26cHvbMc+vqSoFUatTeOz7P1MJao398QEA/EWm9VKLOVcIS5e813+rqK
DfBobBfMGjmww2CbW73vwje9zx60/CSQP0iPqOJktz+wwxHruqV/tUSShj6YnREc
6AooBj1DLjpApT+dk5fVmJMniNLkwu4LP0hmJWw2e3bgtkAvToTCECF76svYfc5u
TGNoIjLWeMugNaFQ9Y1MI8S2YFtnISP4EDNhds9w1Uf//znBYb/lCpM0AoVCEI3c
0deLe2RKv8twi+khKOK6pKR6UUaO34uAtZwawV5jtR/vhR8TBiaj9NzTY3rgh15N
jyUq0D40HLNHSYrPqbfYpVo9JTTRz4KraAz88vjvJz54Xpe4q5AOzBzG57d9z4Pw
8yDwVY3W8vnHBJLWbzYXT5Lrwcje3KbeQoqtzinnKhjQiOHY5x8Cpk5BdR76Xw5+
Bar4+ZEagoBg8ME1EMFkFL6wPchOS0V6DFnA7UbRrUPY5G+l5hSJoqLwuwsYT1cP
RV7lxP7gbwgFS0YkcvWoTRa7ZSvmUe0J6r6WtF+m9dP0/U+mzciBlBl37YYXktqo
+I5YY203lLP4tGwjNy2Q8sptopSXVoK2NS34VrqSaNJF+NElqGZaFXygHLZZoSXd
RZEQX8Qmf5AqYdUAc4utIW1rk2qckBRtNaH9f7+3cvLhMe74m0zwcLDbG1kLqyYv
UfIqkVjEBzH+BL8NGXID0nybMujem0A4VEL8cPc8DnXxvb5bFlIMx4dY8C31In0b
OW02U+FxMJXSq2IxxOKlxdsXSZy7weTmjSFGIgNSb6EMTO8J7RAUc6v8TvAXuNrU
oK9x6dsGcnF1w3slsqhZBKANJMeV8djkL11wIhV2x0jh9p9KI36jJV0dWDhoOSK5
AokPZFP0pP8njBD/PVD1dkTAqTkkBlqfjHC803V5pcajpCUryrMeu7qPp+KHsErx
jEsFz7kEbN6X3BQ+HgALpLPF5sFLXN1wGJqV+NV0ZgaRQEXEGr8vhkcgPEZXoNCV
JjoHkFSyqHjwqU0ZvRcmdyXxR/JlWNZsFg4KM0r4p2tTW18O7IzOIQil4Zt7EpvO
3tJXFjaYDVpVzgwJ55ixakPPgerpFpsoKbPq2gcduy7wfVSndyQ2UCVjkrct5wWn
NZG9NS8gBXN0LCFMIIgLTDGvx8KbHxWGOBWbH3hZqnZVY1shaF1GjNAa0d4WzbAd
sLkQcKSbE3CuUbzPD4QzZwuPTwffMqQfpyTBkU0bjAKqp5Zr+khhtT5+lCex16lK
qcF7wMyc4lKQENt5PO5tT56A9//0fWnpWQl73lrgYWNVIsf4TXHgG2O+OjAV3JDx
/e9HV2H2QrEBi4rQ94Pq+X37o5h9TbTTNeS+9vRqiTaV+LMLluQ8bNfOaxiHlpbG
XYVL8FYfLfq+TKKfi/6nbR+EqP71I5mckCkrJ1Ck2srrx0zVgwYmUxkvJEGEwWKr
qQgoKESD6hpiyPbSsNJ+j+F5RIsppZq86fIgMAV9sDCk63q6x3H/pIPMruWDrHYe
ZC/rjcvP4C/4J0kqT2T3BnPfPS04vXLS9IH5ItOIjzw2b2Y5+xK8G5cjIOBXOuyr
FUxhPkq79xVm8EvXCchmngwK6vnOBC0vhiynQyOcfkIXRveRxm+StRfGYPXSqKIj
PMuPao/Ih9YxLt5Sfb03EgaB3cslPQ48GpwSEVEhCfcPRMVL9xEP+ckJhkV9lhmS
SNsfx6ARybeD2GP+aSxe/ZW/6PCZZmtnzte60zMe6yOdXSDFQg7lgdReCdNCxBXm
pyzSDnoxpKjz5yl88f2QRLzy7ba5Cae6Gpbhp7uDcHLnhtVIttVun3VtiJ0r199Y
Z5HjnSZmFiYgX0pT4vSPQ5hqAom2FnpiZ33yzy+fl+hvIhwggF2UcmjgJ9/qcAg/
H1UqQ9CEs9CmD2obZ22icTK5HvvHMqimwbxgQX+v+/OW83N0k9WfOwNV4NopYqoN
VgxBOi+lYsuPzByOTyWM3Qj0JTkRTOKsQGtTdIMWgcde0ldk7Biz10nsYW3NeYfe
oG+yxMePJAeqAcKH+BKGlQYGYBEr/8WtxZNPUYpMkH24PLOp5dMScq0u0SVhNopU
Jx8ZzOskdGRDL/RRCzEewlAARsLmtOSEwD12l9DTbWmmp7O8diaOR8tjmqCS4ltX
FojKJRIBKnHuafPYmJz/zti7QoEuclXtaZCxNS75IS3/0je2+HX9TWQ+B7YtvNYf
CCPlH2e41+ThTWj3nTmcf2e48OoHXW/OgsXYSmqWdT9TUjuNHFja3/Ler3V0XA2H
w4qaIw/aiLe3ahliVJu6PpcrkUC/83tkar0O2TccW1obfZ+FiDlHlx3xsbeAkpgF
Gt9O7GEPLsWper89O/VG0w5t2v7ZTWfwcNKBTp5h/37/y9fA6H7ov0v1D3dMiQrE
UEZ14Rb80IyuSRlY6VRkQbIIEcsCKJuDRAit3IoGWcx0S6GV59lc1Jn8BWg9dr0d
lhZ9HchWW2+Dsem1vc8ME07aJXrdYSUVI7Q8a0LUM25+6HLAiwL0GDPFsxKTOza4
bsWQF+H9B2lKRkfTrX+fsMFr0L/KVJCDiR77T430AfPCvEccJA+1vqrC7JXr0xHY
a2zYer1JVUdyp2l7XN5WzGnEeXe852d6UOTlaNDjTAAwvjLo/58G/Q6ljyyIXtyJ
F3GjnAdEemoMStALGCFvXRUa2MX5kw3VOtqLwMkzAgcQb9S5mzKcv7eb/2QRAWHM
F51aPR1CmvrdzoXfLbB++lEnCO1I880M9cEB51kEwWoPdwnqEFlO4EtEPPRz1A9y
n4+IinXr0uYhphJkCCP8JWeH0YlEAQVa3ZcpmsTST4dfiIokqv83mpjYpPw0niob
QOGHHpaG+YywHGdS0dvE/93w0pBQpFYJeMsxeSD2aB9Ftf/bdSe+89sBm1nX0Z0E
zVXCSozjE0fi/9eS0ZMJr9hf2ari8JDOrUMkorlW/enaxqeO3zqGlKC3PdzCJecQ
7CMqo1nfhe1KWEAcHaOjgELyCX6hfRibGVgP4iQdkQ1PzC0aMxiFfo24dzUpeBnw
8d7XOSb+/6r26mDOX0c4HMVmNVfQDiLQPwJmdAwiboPCG66T+3yxs4HADYRj309Y
Dg4sVilq4aKxtQ3QDNzZ7l8wcxZ8sHaNEAzprbOAcJdih52/vfQvQ7AT3CfqUU0X
Bm9ErWXbhuS119TtpmDNMVuHAbSGbmY/6qk3dbWvtcfLJeOuO7+gbHmePrBZ8UQv
JlWfnUQTOLeH2oRkxdjUd55kEDR6v5BKh+kpFGJ+kxe/pZk9tjRi8UMhBj3Vktdr
3N+dWqenNEGyMQAWpcXdMdULrOVXTc6vw5W9feX7k9zsIPLwcNeBx26oDM4xRO+n
ZZS8qrqOWJCesng4s/N4rW2hKwhUa9ltqKjw6XROvpWxQDZKMEWaUG0v56DzIYPq
Ku0JgoTgRdsGg/c/vb58UbARMy5e/5gQTDOdBpIO1H0u9K8AvKgouTWBXpv1RkyD
EF+TO+ru4t3xm0QU3xYQo7vNUtbMHjHLalrTCHomYhFU+OVdONwVz1KxLGxTo+us
6EQz21+p2tVmVGoz0f2jPZWbpNYiUhVYvQyo3BKtDLj6om86Q7CLZHe3ziCErhfP
zzvzBqE3tMXbUIvUU56yzEgX+9/1e9yGFDVog5s18Mg7kkMWeNRrzDJMGayWXhCW
wiKpQJx2MGRRAnMrM+zuztpW05JYGN8In2kiIXlC0jc6xS/fj9IVXWUy2Qvc+fja
ITUYjtBApFt+MC+MSgteoppDggGa8HdW+rWl7CPjptHp07oOoxKe1Q8dLrsILLc7
UkBT1x4rJ39Z2S/uhw4z6IVzsKgCrPMNthRplwhuEMwa6Wj8PLosNS/FcIrlTYhz
Y0C2iQL+eB9yaiz4TTUtajd3mdZxgS30xeHl83pvu8YqnJh/3PAQ7FabtWl0hYyR
pnaXvvNlnOf2Ky2agoD+hJ7868AfNeMn4DquzMp/iwR8tCjb2C2ubvx9faHc6vBh
VxXaMZ5dXK11fIsbv8mTptQ6KCEfihfnDfvTkGPsQF9PgbjJk0lW7tUB0Srf3rrF
L5Poj4AOX/Mh0j1aa7n9ZhMsumcYr4QV4DdSNTpZrB0elE+Pp1WGi6HXxJdLBFoR
Uko/4vn/Qi73stmWNBu8Gzvvxlzl9/IsCzSWLVejknYwPJ2kMBclva0YvtS1cbuP
tyBfVfTBtqQUBIvvZnFUSxDhY4lFYlsEG1syBgN7wLpwx/COYbHcTKLDQH2uy/rr
pLZHUwzcm+IGVanIgazdZFQtmIZIg3EGrTdoIJrwOnBmAEkWuXP77ugW8xkLKh89
Ew2PIMcZsqGBbEVbxCTDqDzpogciWhj3S2cYjH49tIEw8eu1rg8TGZeaZvtZjq3L
TF2ZM4ag3itkelZjW7otUnBysiZ4CXTRZjiF2xGoZF266R404/VpSZqOoYRmaHr4
RYB/N2DsDtHAIAsycK3lti0dGemFCUrf3fnCoSVM5y5GDz/aiyxVvk4P694TQhAh
fYo3h3H3G4zpPU1hepacluyuzVsbc/lpwkcKAeRCKscF0Ezbs8RQR46X/0Rh5AH3
vJ6+A5uZvnOJhVHZcmYVDMXJEHuIlii/8G/KaAc2nJQRux8C/NCJTn+s3XsDlaI2
O+Mo4KQzOXOAsyb701wqXeMHyzu67twWdF09L6WYQqFWtRH2aJK7egEsQpKjnVoM
HdDzOvSLVMIX3/W84lqzGx6Nf70HXpvZ0axRpfi9B/lqEfn8bVbGUzaI3uf+NNfd
VnMO8EbuAwysPhx+BglhIisQyhVS/a9aWrMc5Ra04sRJFq2WWCxwQjfTjzclvWZH
f4rASC71SJLsVruntRk96PoL68F1EoU3UJZyP5JPYTxqjOFRNa60DEfOLkiV9OFl
6Xuhdn+HaJxmD4NPR42ExvCRM7EFujk+42SIc6r7x1xidJ08yp9YTFv0GZe5nQDb
qooN33ur/UsmG8bDtbOCC60AY27o6pLo0vernTMWzZ9h48uV81kZpaMUfzK8xFKY
w5lKmuvA0COqtivMvdNqMR3uXymmBXTE4eGJektve2CErBb4S0wdgfXlVpo9dwFT
+iaWwLRERtsc8WWDPj2iv+3YCbYBosGwOLqbuQkFQjuwPme7GsIsZzxmyAH9DkTW
2Ec5iTvPoIlGddbqQlIW8hLsB/TphOTibHTnGeBx6sAq6zIlYoaF7h3q5bUKQ8ge
VnAKSjvcy3StdcZpXALMaUy6dwYJTk+eFpkJuKXQOKX8mjJhbvvwdQ0A4N+5vAe4
nZnMXx7XpWJ8jpcH0r+hVnaAXBMaQKsEVVXBXBMI5b2V83dJYhv4Wm3G0ctjK/JS
NOPvRznrtWVGRWQSEuKG4gRQPZXNut0vqu0z9Rfbc00PqmAEtdLExfJUWi30BQ9r
eL2eDipN9SyBxPewCwYywIdB7XP5A0QBv3boVC4EU0/b54/bsB+EqdPez5jkTpd9
SxdB/tNQcMRmBMRg1dtUDssKDUx2vaVWx0BbJlDNrzucDt4YWUW0V+JahA85LlMf
fdwyocrqIx8Y/DCp/BANyyL+1GDOTDroR7mA8LNvhiPgIrxcnWtVYqlRx8aNqxc1
D3yyajVKtcdqIuEOsXvW1HBvWGo/V0cUd7bbLZT8x9ezQr0mUJqVnrMu+d+Azw0+
uCuZXmdbRO3ObAhE1BC0x0xN1qx3sO3Nf6ptfKbhWjpWI+kRLS0ayqY+DbS0y9cL
9JCk8pk42SRml6JwGS0+wvtyN3samAQha5ScGVvj1x/AsH2/lF0J+6GAnLllrQJU
lSoYjA7gdi3sbnB5KlcUI7qqQkDeDd9VpM/UOOL81vJGjwEUNYeJxKlireVN0uOO
r/Vbk/TjsoGxt71shapoLjd4JXWAor1sOkPpXRLlyk6GG7JOVsKl7Bpy26ECS6zT
bDvJJuRHzEcTzBsBeGhGNsiEJaws4qUtdkJJO8AvpUyjWmt6mxFmqNYMfd63JUgU
pJ9qrTAQbhVdQOg3vMJ4z+WhQqRS4DkEhJ9vycfIqRBk/RzZgMrPJSx81dbyC+US
xVTyvlAzB4LET5v9VCpt+b+mlPL09VTH/pl2ehIa9c+cwRK3Z8I0krP1tpqZnRlD
4NvA5IUdPaI9Rn1xBAUKrxuG527Tr+gXITjLdt65iG+G8aQ0vPjdM24Rp1Yn2MWc
pEkVIAXwDoBCnfgiHYxdekteprhj/xSl18iYAHMCoJvrd+GktT7S9XtkIK+7hTFB
6GzgwFuvea2OtAio0Hu71XIAj/HonjZqxjsZDx9MVr+MWaKqAzq+EJj0m0HWzKf4
Dd7CbyAND9cUjeH9fxOYAMZyDqAqV/CocwARi2JnJ381qaKg87v77s7vDNLhvTF2
ppPcAgIB25NAwLJsp8vjMJM0I3EdUUYt143NjvrAGOFIhfoPcOaRAZR3qR+UJwZH
EOiymwYnSsGIekJza4zIylOeF/Ufz+3HUuek59ZXhAi7Bi3WjyttoQqUr1IzA0yT
0oD6xSAmLRuKs8sWc5N3mv82q06buVrRCWGcTjDrbyTvY/ymLvjuGD8gsVIQALX/
YJpXCfH5w39eAkUlFfTEhyxzTIZuKcH0Ny5ii7iZ9vgHJrnIycgOAUSKLOkqNDij
XlkubuNjqq3sz7cq4KC5z2B/RUnMCCdlCtlgDnaZY1WCevlF/oVQnQIbp7T7WDdN
vnaEplOKuE3PQQDr685oqR4aWE3A0K/qFx7RWF9YI4elB1cVTSZ3LVuvwawVdVq4
OWjeiVU5ZYVZkHeUFgl4sfCVQGg4lLmADceTwqz7oJzrYvKC5Abmpj+xxo6GQidR
BEdq6qSuxF9ONpF+A9rufC0CyQUkNP0CtDdOr6S8LPw+Mr1+BMJa5ApoH1o99/CD
6oy+asQa/vK7CpVlM4gHWUmON7QY/qjSqEaS017U+japgdHNPzw69UBFyRDQxaGd
eDu6xhva22BXoiMMwBUWyKMa0YQ2QBHd7DnGj7+ogK3F9A8S1AWjOUaK+YPXeQfr
/fpKiMPKFq+JoamMVYO0p5ul2QEZNwN0klTLBn6hXXEl2pvaPiCGfNU+7VHwxgKA
EbDAr243h5OducX8hN0qxTcMh87rMMWGMCTLygSEoRazG2wBoVlyyiR26GZylhb0
CtU8RObPxAxeyFjRG42XP8IJ8RfdHFCgU5mpug2g/pT9FTWEdlK5AJgZ2lsLWHQS
4RFuGxwEsN3dVjSJN4U/4ZGdWDJGmyJuGL3zpfWLRqaMfoggxIEM0A9hOzuNH3BY
xNUYHSEvKSEvEYqyI8iN2nJZ3xKsv2D+ux4DCPWZ+BwZI2hpFvghigf0rdhoUE8o
4NCF1C9AngYLS4Sc9aO4VmplMv33oVH3rojeIm+GN26P+GgojAI3QCHwpC4O9UTP
aMMW82hZspQMh+qa6w+Drm2Sf49iiDUkvacSHsKTPLSuI5V1gqz2/vyvf+HCYMHd
OQysH+5PYog/IiRAZNSLL9HfM7LiO5ShSOz4QyvHOxnptwzp4+QDl5hriR0oPVJA
11IglqjD0iO/5zzmDCBZ2hcEwp17VpPOpI4VNfwuyTQHJGvABu3u5VXZQ1F9p1Nd
1kopTQCsjYr9CZCcYBfzvgjkpBja8mv1LeNpk+A/1p2IJC6P7hrdZazHkgS1lncW
o271bXCSRRteBq5LutNYNe8G3p7euuVPRajaNwghmo1DFyNY1s48nudK5TdQm7+e
ChUhHI1/V00XnQsnTv04pi7oPDYbHtfDCkbLOKfGbPyRu/NNbug+YzXqryn6nyUY
KpHPoSiUcyh62Vge3kUvEpaUpj/V3cxCfzipuljRBcCTYxs+Jdl/g6SasdvDEOz2
cVXLy3U9/WeHF/aEZGBfIoYhod7qWVSKXI2n4X+PxmTAXTB5HF6b0CorEiaMunlt
YXom8tDYgT5xcCu2AKLTegfm8sIutXIacdhW7vArgEsWeeqXOslC+pqsyWZx/Bwt
lClnuBjS1YjiccEKCLrkBVwlZqI9kTwobbLLGAhdbKvYJ6zljuYE/0c2yWbTSzT3
zro3oGx81eqdZ8adNOt6da7GUdzdcUuu3FzpLPFy904ph4/IKzoiT34V/P0Ep2Ov
Zc7YXkkjLYzs0xgwfJ6Y6HxUeUyZwIaFdiaOSsvTobuDcHS+bTuPZ5yScN44bQrC
RiYFBa796Z+SJkomykGe+slB/esHPPgQ9r53SIJmP1dBN7QawMkmrZSSq1aB7uM3
KrK6dxCK70VkhGZsKiWfkR5tMUdyUrR0URi5ZI6bWyocNv8b2uC+JCIBnJSgdOmc
RIqV2CxQODJv3EikImOjmu9QctbBbCDQiAVeaUoNa+iRADzyjx8KqGE2rkwR30kZ
j4/9Xiz8QhboBWflJrePySaRe/+KHA/IdlTVsMjKKQTEEhrJvHxXx2EJJdsJ2wQ1
lY1HaVwbek1lC7vDNdizBogmyOZC4qoxlrFYzsiTBoyQ1yrgrVURc8v4VsD8TkCY
viHmtGehub2DgIEkHCVtjEKaFzISvRGM3AUIwB6VO36xFkk2IL1IA+x1+db6mv/W
gwJSMsU86HkI04ZXcQ839GPArO1R/sDsrnW8mgj4yeJsQH955dpSj7yZagRJjAxa
RLHkCA/E0i/6QnTY63PUHpR8QZsX58JHHAiNAjZ7rJteNNGJPAg9II5WQwCu5EjZ
fUzRY1qVSuj4t0+VREGlw+qRXr93uXSQsPmlB8hhh08P1GF4EaQXsVQcN+z/dyXu
nkkdpOtTYKvEMrBz7qYGETe8xXcjVAgtTnG/iRv61sJJ3+jEl0S+Hgfs3LGKGq6L
7d7qjo6OTgr6RVGesiAhXRUGs5PVuJUGAnNcgTWwzdOL8gP3oAuJlOBRqRFZtLse
keGfNLYLhNEOmNPETXFCbh11SQlqaqYL1eD7tnoPvJVSevXL0YlUC8cKUid+lF36
GUe3BuuWvuNfCR/hZhIMYNIyzuFYtWGNseJvSJTJczsRBQidrHwl/CCs9BfEvNQg
0oDd61CzY1vepYBOKk2QMMgEGpGocuowxyD76oGhOtVS38OLwpNyvj2jJDGulRDL
trCR1uk1y8Cx1GDf+xhfo99XthsnfoNFqTGwIZtSB6o8vWsIZvVty3QZDIFOzsbp
CEV2KIXVZWjAPPNMtPPytq5BV79XJ6rLvv3anb3PI5dhBLXSQBSqxizGM80xv2O9
lc+fYc3HMDL4oEnbxh9Oxg3ntkyRZmR2jKTRhLCGh92XjwMWZIdc+4ZfqhJzIjoK
npmtQCw9mrbQYIC1IFWC+bHS9ZI6mg7AGcmVEKw3owPweAanPguQiSlao7lQgZgQ
8AakT8GL3CU907r+Chky7W7ecP56y9hfhrD4fZ8kbzOe6E5IR+X7v1qYdwTLzChQ
U0nKOt6SdiTCOFNuJ+K9J/tbkdJSkYNnoO//W0yG6BBTGT/AQi3tlrzizM/WlRcd
qpk8nb+WwfELa2OGG1GoVCnlTpcVM25s4QnCsBugbd3hZNzdq6JvzkHJd5PAYuhh
lStYF6/F0BcXYjzNnrwI5LZDGakSfhXhDViAuHJUZVNBk/u5AVOHW1YrMwYCpyba
fHMws59LVdKJLSgEwJSJG31FW6Cu+cePOdSz0xlj0RO3dfNGsibEB4q+Qy6rnkE7
EFUDhVkfl3eh6CWbqVs5FdHtlDOhq2lAhQRtONxJo0g5lTB0mhZt6Fh/Uod40Sqb
omJtJQUuSnBQsx55jvv/50GTzvuXGnv9p7H1PNmAKdjsWOoRAiCb5UIFYtTOzTC4
MbQm+z9ARUhZtyevOB0q4BnrMzWJUGEt+KmNFNi+mQ+DBM0z1Ib8wiCNfjmPJ/kp
E6WJzEJfIFEVAkfQuKVVSrlGPw6OP/x5/nc5M/51MpjNcBIOoAH868Yrel+3UG/8
cAKICkLnvpOFVu7A7vuq3eC9sPwNp6uBJPl5ducHaQ6WN7BJIC2XOVBtXCbqC/kq
hI2QEijAHZ5+UiMqjzim8p+jU2jhyG7CHR6LZ0AhS/7oAOBkhvCxoxq9mEZDB4cg
GAeWEtQTZeY4aPjrgrOR+r3TTE6d3iYFvh1hckPw7aiI/+jNwCwp9buKRVgDeeXr
hSixfpJpEXrhvk81yIp6j11VYh83f5Unimzoy89inWf3YHPnMa2qMV1xlVeYGS7S
SjDpzI6PjV1X/ES5AeWp/EsEvlbBXmG4MUM9N6TSRYXBZnGntG9ycFyKmXhHVIYt
/n14i7xPUpN5HVvEpuvzkMdxEnbv9PpybWmlwxK7w1Zx/Xhj2owg1dr2Sz/YAOdp
AXzwyQf5zX8kndWYC9WohTZMIVg8lQoLf4KKiielRYqQCxKTTO3SJ30MlIDRsfui
2Az7EpFDIraqWgKKZ3i74kULsneGnfVoezb2Z6WSUf7KOaLgFbO9H7iavTwIu3Mx
R5JdbpwpyeXmK/b/8wa9Y/orPoh7pBA2+dp7s5abNVnrWYN6opf6TcHN7FZqjIaL
/v29syIehZzq8/wyeLJvqQAASWnz01bxMQps3jJhO5iL3mwGoU560Ju1bKdY+Xbx
OJI9rT+OELq87+VYcwYNh/s/FgYN+PGUOJHqkrHF5qbYFPX68jKNvIqmRqs1Ept7
Yn4tzkGUIIDV+MjS7e40RmKu+SJgJgBEcbP627lkFvtd58Q7G+NvPrMGOSjtlCyg
lHQatoZThnYLhAMCfWSBhaZfd50iJvKnazwBSnrgYlCXIKt7UzuZNUFHIuWbkOPc
bq7Gy5Dx/96pGpDV7wQIjeAoTGQ8DLXiFKhSMnqVWIUGaMtw1w30vDqHDMZxuzPf
13rmzcUK0CJIojqdeEGamaNipQpeQcTP6AN9qo+cyiG7y7kGs+2uGhTi8YCQl2HC
X8ZCxYj8mP40mDlS5h7J2Q19DXFXxVSpvWigua2nnIORi8Yahivh8BxIe7iEi/ow
cmjqhAk8jcs+2Hpx3DaC9Kyz9RlAM9MFLktj7qp5RyuJLW8mCQFsXgeglVWw8BJf
r7nQUuWudb5yxIO1tPqBSkthttz/c5dfNLDrWcJw6Uf66t1Vb8M/Kr38Wu7QwPzM
YFC6ExG5hHnrVm+cttJE7wrcyE9PnbSALwyHR3o5kXAodEDWVVKfHaQZIDJxo2C6
oywlh6wqg5y/7rxkCfCDPhvNcats5obn0VHBghaFpq64N6bLdtMr6K/1J2uHN3FR
ivP+UImmFvzwIrwA1O9I5yT7sCXNnfKF9n4MJHHbM1MjzG4oKjZcNSNR7IrWXbY3
oI/d379NczQ32nFkt/UwKk2QzZNhqrQIn6oUWmm902NOS5F1t4S9y+vLsubQG+YU
GXOfIC/evdRBEvKOq9mQ6TMA2fA5A/+jm7nnkkK3JzTpoc9tIA7FrVDNRa5Gp+7L
W4YegyCJMF9eyd7oJlCn4I/Uag5SViNcUkDhLhkBFIJeVG0Aggf5RtqGtzO8n0Uv
xTroaeeSzHtRaHv1O4nZUrxR2tbsG6QaC5VhsUi4sYa/41H28xxpBzwmzoUHow/S
zympy8qEfH9LX+qOW9JqqMGzz5+t9/zjzBuCn1MQiUaMnL6ydWeXO5OBsb5enGMe
iGw+Fc+WUeMnst9bymW/61sBy+2ZFuxJWrgLGvL8MFJifF5QV2j5+KuEr6JBiUvs
kLYuGv7M8l/xK6EtNN9yBJyWec2W8GFDrMLXQOJIbRUf8VJbJexdViUlHETgLIap
I0W4jT8ihA/xLrGya1JFUomb2U3R7xzjcImvIXqJMv3Uxw8l+pS6uPwrQr/WKPeT
qEb+HQWgZT5+eYHE8FFLT9JE0iy7Jl5qWwkVC3bDl3/0bWcMfR+0OVb0fC/wi2rL
Ia9pv7CXnxkiKjwsgVb6i4Hrj7bWLxeT2nduP5HDxhVq74TzScw/6iXL16UDpv1a
CQURJE0sxG1Zbo9Givb/JrH7LBUOzHvHEFVW+KsH2IAN9jImNADUDcVW+S3nTj9c
hzuOCUQBmHBtoHwBuyKjlmpZpIbtKYvs5WgWNMk/M/XYKWcEUk9HlB1WHZyDnppC
bg3huGOqGlzlzLzBDR3udCX/eo3S1WqBQkiNVLQ39ePH1TioYN4f0Tsfh6p7KVBz
JhynRhovd9TOZgwZ7tYoRnrrAVcXIn49qkHmbY4CI7FqUG4UBrd1A4jvKuEqRq0y
3YvbBi8xBhJhIANwTLCSQVwS3MndGqomkMaqz14OjBDoaUvhwU1u6TdxYy048Cbc
U3Lh5dHT4XqNHXw7Qexy8KdwCGDCsOtCJXkf5dSS0THl5eJkI0GeMgA45U7+srFC
bl7Rbzwunb6fUEphMYuAahPuVJV3hoDB/cOsZofyabEZ3oA5UqdUzF3pzdSagvsK
PbSWWKGWVFtg6STlHJIgitj+/KSIDnyYOUgSFikql0BOLsbH1B4xiIr0/zQ0S6GR
HzTKOUb7AtlvdlGRAn8TlfMCCLrtzb3llc8FYGRV0ufsuMfjeRuH1RpYd3BfXc6p
iIn83BIhahtnzIhDBkwaU+TJFXCYeRijoK1w8KkVxlfPqI5LpfX02iXBJprJ5e0a
gfJlkVB/YFYaKIPIUkv2ab7uAvOSXAJ1yn2QxmL0PKk5C55aGe9QihD4BP/xx4cD
kjQ12Tu0RAu+QhGGWT/r8ASQY4+RQf2XLu2Ls+esWz0MfjYdCoNQCXSH6VGU1vKD
dmKdKj5cl86jpE1Vesd3hFUOlV4w/VERMyal+RBBUu5CJgbjI7dNg8x8MlTGgueJ
dwTnaEouygYwqG8IFRppyhB8iTgKpdcdjzG0+C8IEGzG7zVO7HHTqXq1Cj+ParRj
6kdqN/PU3O0fuDp5BM8g1o6u5uDm/bowlx9W6uzpDiojd7JAnDlEcTCxDmW/v5GG
eY1PDP8+LBopxpuOLWfUPDfNxNzCY4ursusgfZx/Okntjp8zanzrn+h8jW4vKceT
mR9wRafB2hbazN44x3GINcyP9eEE4yuohdQ6IAJCAphYzeWN+dd5PyNJ+AW3sNyC
Rv7N5Qc7q00+rXWfbMU+M4p0DsaFynEx2PS0yBKZWPIzmgA7wS49u4Iq7pB4NawZ
zVNmA12ZZgYSCcqZYf9QyXFdSVzbVKvaceln7UQaVcBjaElm7ydE7L5Et9YjncDo
M+nX0ApX3H3gbDtjK6JpstOsNlGu7ZyqQ26A+lw4azrGlJCv12jTBD7J9EJe9u7F
/2vsHEkDd2N41hpSaqA+/G87R3TJ1mPBYyiZUs2vkdpdRVIuqpS5WxEJq8+97/+s
MkOF2X7IvOWM76yc3DZ1wHCWKE38Ls0CiVbjqGllLtt7l7ZfGEIWnjs7XhtyMexg
m5GvGnxeXm7saPVGJY6gVoAYhKIRS1k3DaNUXBGh1+SeB6kAYkIv0dxv2JglUKwf
aPxm7Hbt73gJl7q+SXPGpO75cpr27Kt1O8K/ecpo6KCvUpu+aYK2Sb2i2iQuFgbC
bbpSo8uoXgohwMjGfMqyvOqVpOIulQsiCXAm1kX89vt6XijvFUvFFsxNBxKTsDJm
IDDOOvTQCciy9za0NPlOBDbR0PqUMCukU66ev3UxPeEzFIY/MPgd0eulBTltfsh6
aU3BYekEv2B1/SalP+d5rUu1JavO6vFys3mPX0ti3SRJjDbboV+pga/HkYkPxN4v
AZVwUJhnkA2GZEoKPSkZVYfOos1/nbLlpDpli3KNzU4IpKPCtRfI3r/aFjx2aGQZ
Uu9RO2BK2rGFo7Y88F2WjhBEQLEwKfgm+8V5RvTCkGSC/8okQBqegOOKyuxqCefr
emfvvVkQVbxSo1OyK15wbKr7Xw/KC+JcNGVL58PBuSUEfdMfz1/wRmj1P9M3aL34
72fNE1UqfigyUT0+6dZqZSAy8OFF+VSY8hvlL4HZpRNpAK8yCG1GFEt78LKYvHBN
DX+CefHSw+hk85WRM6bI1QqkjykCAawXt6+eGaUFlCiKD4BGuq4gH3E96igE5vh1
W175YOyGKT/UfjPxgVe7696JI1SRivxsrPQFsormnk2qJVtESNPheXuji0AjbVBz
uIgxKpHZSMUqXnDvLvhHqQJYO9qautvRnUNFxQVMcfIPdnJj71Zm464ITarMH2bw
8dw8Rd8Ic0F5p1rRr8dQei00EAuHV0U+f9X0/f9mu8Lsot8wsm8xz2hvxKF3lWd6
4cRmriTI5xYiwPZXTwBWU4Bxqjv5rCFSfwjorZ5Asw4mDEZZXexcyo8FZ6QxtrPJ
16KC0K4yq35k/zvbaClVV83JBlL91ZxuExd3oWG6l6RnRUrSZhZ7m0vHJXJlBiYw
5weNtcJ4jk0XTv9BpsfbyVqOQVyyS8BokVv13v9v0dU6BBTS/baJjXKni5XawqqQ
R0eZkO4fu33Xv1gNhPjTnTZjv+zkrN7gLK8Y0dDcf5glxa++eHTzrkAXA9wNDWR4
ivAlvHvkgGm/0UmH2mfh6oajzd3ToORUGsE82AU2qid97nsFaNqc2A9pL149QPfG
q6uE7/o84/lvunyJANSn0IRssN3EWopkuu890CiCWEj9/tDdGxNS0iydZ3D3gP7H
Aayc/X0kIDdQphI6rC+nCG3Gh1ZkK+JYNWMRTy+PxvE9P1QCSse/5AtmxK2rC6DC
BVeVQAPjtbXIjyOzxScs26ryAoUWuBYTvjFr2gMZaxP6cATYFPYRyaLmymkEFatT
Su5xNnzmm1MHy5gtIr+ZJEaARdF/ImEFv15bf2oYHk4XQ1oKNsY76SafPeKnsQE7
wT06Gw+a2f8vF2AslNmzi+7/hNMkSu4AbqLOpwiRHiR+JzPVbGTwRTO61N2+g1Gd
90bEQnRZbj2dnQwclkXo9++7W7vfnXoHiEomdrhakeLqkBIPeyVjSfREcmE7FxeR
Cy8RvaTeKBF+pCIgJ+JJQ9Tg/Z7uzMKP6uNlK3NCoRLhCtdS2CS/fwnKKuwD1mkM
YNiANGWIjmy3FKW5kzFDS4xILieiluMqgGZXahXUdeIxVjOnTAj0O4j8caZk34iw
rTTBtf2eBLrmvgEt99TUbe4BociWUhM6n78fhbFa8MiML9tEUfric8ixCv8Z1Q6z
I9ZWfmrnrFa9LFf3RnIzDBzveR7vaVu0BgxWKIp1x3iK4jeHJM02SIGzppeVglOa
6/KHGPbEgfD4PPTO4raFDtU3359a27K5k+z8M+jnQLZrZ1UqYB6TL6M9wpBkvbgg
/Ax0CfMAa45guiOqhEDGcyRiG5YvhpFxLybRnqH/b19rewyPEOc0zkPwM2TWohWK
xt7i1Aek0ZLQ339HzusBF0R+Zw25HSjeEfxxbRrjU1NwA2cr5Qilvb9GoqA9+eGQ
jLOFH7dRwqHOTvthHZpuSYrQaqEhLmrtc05EjxMJ8pwfoUCi9dXYtI0BWwUd72DF
UvYoGM1sNxjm3Xbe2Z2IIIxwx1rSnQiNbJ6QO/j7Tuk280VuctW29xB16urx9iFz
hku3RJdCnSlk/Zn73h9FqnyMTJl0PnuCXQF1t+yD+CCWNsMvucIoRmArg1voPl48
Qtn27ZaVMNRXtLU9c/ZDuQxjJNiBV2Z7bwbkGORh6onBSdeiNg1pk17hEoUaw4zq
n76bYgjmCUdgOobZ8UVuaIbr0FRXDJGjQ9p3QmS3DoKMIqj7TZ2VTBENHA7EcO9B
9Zt3ApmdHYWV2yIz3M55xn/Kq81os1mes1qsS7Q0bkh2uQaDfehQZTaEz4Cb6g3n
Q05H7U+duxUzlEUMipVx6Ht1cfujZ4JJQSXlpO2uz8BEtjsQZj2Cg9atcCGpRDCC
xhKPGtjY6KDhGOYENwLs2gI3H/vhUC8/BMpyw950cZA1CWaq1/qcJdMMp7agisww
HnQrIa5ckZSDW/9EiEhJ4qEaR6hapMyJKYSA7Uz0g8+Cee4lrqZfNjztB/5YMfkp
Htacm+Vq6TaOxW5VLnashCEVqdy7QimuHXrmaX9tAUQcefuS8EjMjYqaqzVW621x
DqhW65NWcWtuGYVRLVhYmq0Tp335QQPRa0PS39Jyg9RRQwZRXwRD2B/Rh78laI+e
SaaqHfj/mVRGoT26dLhiGUOjR5QgeVipPnBp45E8mnErMfBvUmdcHx3mnpX79JiT
n1b/KfZFTWIPqUXJzQBp4Xh+GTX35MXy3OB0UF6NnnPL0hpqIzn2lcqN6mtR1zJZ
EWRIxUPj5iagFzyj1tW1i/ZWucnye+FELG03pGSkX0i0POPGbm1BbvO2Uj8zAwI3
qkF8HY8jalu93jlge8czzJWTQVnAa2Lah2yMR7jN1VLRLuDmY+5vlzDvSghjGRwW
CtLmoLf9NbnQK7tFzSAqeQW069szPYvkwT85CrbsB/Zv2A9DK0fj7wdu4tEPRxUR
eDt53QpBru5b5Mgk2Afv/w0gIeacsM9wc9noTWIaO1ySqBlLGsjo4IDM2RtDp+8p
BURb4XSCxeIdG47DYzpuRHEQwmKpWk+lPUb9mthn4TvkcOr/WHWpqrX6HDXsuTOy
MvfSwrmnUcFbKNyOl35qKanoAM9x79rBcrf+r5jEgmne2TEL2GUF7bp1eMMUXLQN
+TR460SpxV6Y7UEyR5jlasuimdDydD5PV8N3V0wkj6EUZ6R7AuEvxuWtW7qKR9jD
DSTTbYzj8uW0IiPcCkUSntDJUUWN7TDDvAv4vs2duPjcC6GyR7bL4QFNVqg3u23t
fqrUB0vA+O+4n5WVC8JVOdD2QrnDw2gYc5svjVbrten3LmI8ShCeY84vFgM2KagO
fXt3qp5QSLr/CVPit21Qt10DOZIuLL3ZF3xL6q/nYXF+72uiqAgEP0hmPO5uIH6F
FTdHYcRWzYAGeXbKDKLsY0HnWH8WpLuS8PLv7DPUNwkNYIHMBowp6e8XzX09VXCN
nqMluKc3psogBK/N8P2aS4JYC5bT9g0cG6gBnvQ/QSJC/9yiWOf7/R7Jaybf21dA
CodO6X7PTTB31tD7jq8IUAFiIyXGO8qs0R/yx1S/6+D1mz2glkYJjhtOkf1v5/ht
YOeFXM3QelBbeENOn5oOGR+GhQ+3qoL3eNGyuO5u3kEDD+0DS5bfRwAC/L9rwyY6
hVHMSjiVEGn0LwZFYRXTvrYjauC3etjjWaCCfRlEAWpZuTYuXVySiIH8/QR5tSTF
CbKrsvcmLkZqucQakyL91VOwd90AbxxWexsr4/4KGNMwQ10i9gyo8CVfAL4LHYaH
KO7LjEpayL5GrATUniZ1kf1nQZldr3bYQigPiiW6L/bmnqbZFIAwMG++iksGveO4
ibFNVn31WnL9mMQcc24ksfsD1VgjFqjeszx0Rg0mAwgSnU4CdHoLRXwDJ7TzBgmI
COXxB0bkY8MjZ8Dx4CL3LNe4GupUHLCQYzq4ghGOgCLIJAl5Z5szsCNiZKZeCpEv
eU3WMdBlwoSzIgdj0tB+9bvGmjDC4YnRhhCx2Nspt5HpbPISXxBcR+BBQSmgvsBA
FQmZ3zQbKYnMaLMCyb2eJ+YJnrk/LcNfSCIrMS6lOgHY4E+WQ1PBuR+6MFZqMc1E
zOvA9B+Vl+MVtZ0UMsbv4BD46Oql0jk/t6h6i/Kw/umWDexSiiaBV2U2Bue+4UR4
ccXlxwPR/+Kw1rzObnxvTB/wTBxz64qWN2FB3P0KlYsJM9MKlw1QpBTK1r3Lv71G
t/Wo1LJ+HUH99ZXqmITLytCpp0WLYV7uRESzFeb2o9hmD/Y6kBn+n7bLrePzBhR+
8kJvuSrR11Az2vvzmuTBcOxXKHksiuq4R2ku//ei3E1gSG8TAS3qMWSKk8NlcWnq
DhFJ7OMkcwf/FPm8uCO4BIZudQ3fAXw7hq6Ts1q754eyVnsgNtpwWBPgUjRubDSI
h+U8QayBSTLKkDsAtUHbgJILzQs6Y8e39gJZYy/jsbbhgzuK9QwcU74iYW9/q373
OCB/UpKGG+zTraXDeCbwf91JQTry4wsBcpCf7grZxB19o0NQ2ZMTv14nMLvTVyrW
LS2L8ZzbQEgbNTEeH4vnQ224ZIZq0tkAKmbuk/Py1H0mCP4BZAaB1c2Gp5KBU9B7
9C3YfHppaiW8KjA/f7Uw1OmdNeyCXf16hyiakSKICMVr/hGeaZL9f85djiNzMPhW
xJbDSLAO3y5m5cyrrcWd3f7MZ41UQ03A4u+6D39NWoVIIBZ7VuKCgth7NCTBoLLD
33zkYRvMHGObjGdx/6+aFAWQ+gy2maCH9nbYpyWNFiNYLBZg1BFSkOAuQAK1NcFW
392qcOUHk53uZD8XB38qjXkHtOFOlzLaXYZM7VUeWl8JceX1F+Xawnm9iH6zBlQ4
qp8tItEiYqdrgaqVxCby4HgLBWaX7a1yNk6BANe7AerxlN5A9ZKn4uWV5wHo0Esa
jbmo/Z5rkiv96N3S7ICEfxigQrMjwlO8WOLvhifC3XimGf+s4evfF1zUDR24UX2O
gMTDsr3tjkvxkt6m94YJH9GDppBbcmJDukvdSp7qxXVgfOUeoZRcvuRoaSG5yXxk
pBi8tsQR4riLj3zmH7W5Czu+jBXM1vwhhUfweTFJ0z/lM97NzxogkaDZRbNz0UOQ
3LUbtFc2gkHc8bTWN1sRdeVFtIXap2ys/yBcmkTU4CogcVtp/DlYaScBIoH/QhSU
IniGagvRP201yjNYhXcL7tRh6GcgWFB9pBCIMTQc4OzksMW0taw8kcK/OVEEFPC9
BS2jQqiKKO4RaqiSq4nU2I9dtpNRtXd9lEkCnIY5MNdoVv7ZSK+w19jmaWpDP3gh
R9NYhVqcYFzcomqT37MuxamG81NBDAzzYRBaDbrd4w2wRF9qlmX6lCgwLaVMVXfT
9QQ2qiCS8AsO8R+xb9AJzUySwymOmdlDqcf99CTdn2+RhScAsaZXfQQZbaMGXNSi
3d6NdIjVes1AaaoFTdco3vesIPquwEw8GTX4S4Gdb6GKizBpj3w3a/XWOtE7FGdS
RKoFN7pKRoufy4U7jSRWIspZ6SiKEiKelZFGFBCWgf/nZcjuIqL7aSPctjynrXMu
fTBcj+qSCFe5xGI0sb45DHij/K4XH1htp6p2wDlg8sc/HJLFlLk7sL2GqO7jxBcN
q6JbchxsEURioeOK8HqmVzot76U1bY2kpVQH0jtSbsmeBJbynpD2QwbbXJf9nss8
mWUmy7oeg6S/9mJ8ysYuSGUukUDK1RVYDVggBhaIqxCFJ4V3advXOkPm+/qCfXEv
Q6zIjSR5ILJngFMjRx7kQACLD8jfLTNJBRWSKr97l3WJrXL7VT/gWIkOUT4AzYaH
C3V2dBay1v1aZDgRuLrdfow3nknnhaK6oMAS7JTHFDw9p9WAE0Vd3WqfyIYLIW9q
LNgeZWVnwmCCUKHakpMCgn4E0fP4v1FHveLnAbGbseLEXUeVK+gJAV7WdRUQeyH1
IKArPHLYUtU3U/1xhYGK0O3ncKIOdV2MTkaxp6iv0qvXrhPgzmwGJb6hvLriJyNu
Sc0icDu350t1m9NJTaWpMI9Tp+kln5IPt8a4X2M0/5gaPYAiA+VEjoQrlf55WpgN
wVanueSlV3KBKvobUeGGp6ju3BCM4ltbk+6Lz6hPnEJLGWSMn/kLTbVO4GVZtlfH
BN3wyTMrx6MUbdNx7XMAALPow3NXVzzOWvTMYlWUogIidvSoXqwnwkWcgUGmrCaZ
M3UfSfrpx1qDHFxPfw8/1hgiYEzClle7YOQt2U5SRm9V3fOMQAdv12+P0IkzWUJ/
n2dGKJ/iBqwKHgZ0iTaW05LT75S/0/lplbtICJq9NP1HfGVBxfsol0kJKMJMgOIk
5/4WlFkyeTjFSbcJowWDUS+BBFL2XD/nq9eNAAPvsGpyDhRDp/S5M027poIK/1UQ
JSFFgGQmCvcOYwRyQYrU734lhD5UiYoaUP0fTzpHxOd01Riy/N9FaXCofCPIvlUb
19NV05zFPmDkUePQIqgunPJLDubsR9nFLRhAq4yn3fweM7wwUQ39r/JZ/m5UeLYP
sqoqt7mPBfN5GvBD5bFBh/4ShkgPEXWlajn8Z9KRtknvMgw/88mxiOebsbxVMP7U
kN0pfXf1RV1ke+bQRBDPgaRjMAnjkRmZNFBu4nBDf9oeH6WhoBn/Anzp/fYlKEmF
55nNs7GEd++0wBE2v7lO2p4EeCqY2R3CXWUnejXlsqRzvawl4q4aNYnNTvnDbkQY
Vzh9O3ux9yZJGHJSUSiIbk18N6si8WbLrv9bKzj3t3BWzeyYNVlt5VJxPRAdUWn3
6ZD9QjNnpPV7sYGvSPmcYi8LE5XxbPE4pGvhF5lVEpMjSdvv/p1y0+y/YHpbW8X8
uABLkTjkfe3rTHzYWzq1Op94B7EatTb9UgmjdGmff9114lDHud4UPizBIMQ7PhfS
2Q8Bz48AuJ8I5WRdsa0o5OVKeyw2rmDSxikPvXPGWnrUsfYfDZf4vvb/KxjS3u3z
Yi0KfNxj2qbzQxW0wkOJ72tqm2HmskKqJTsgf9+58vaGfjn5Vo9a3pC6c1vwhyMF
SObSnQdwpaWsdDI6cSmJLyh0oiQ9V8puDZhI8Wnd/SBP3hxIj557W488zL/3xTgI
E/pOcfrRPIgiLoDPBlDQWWBoDaCxEdqEX61wP2qSTc5VCpTweTsUeC2VxCZAZnYw
27NM7q+ajyOpXBMwFOy6QqybL18+YRQLsCk4dAh/B8a6KMsJdsMhJsNh6Zkdea+p
lZkL9OyHMzRJGWht6Dc93AfL38i/2d7T/sUu68BquumK+8XMFTdrUnelGtRDmrdv
dQAoGKT21KFT4LGbfsRWhkNHRy3zzt2WfazZSX/+kPm/3/jHgceeushlMcOCXsK4
z8bH5si6fAyxZGjRGvWpUyCyaRe3Ed+AVM109FyUFkeJWYEsFPq5Ld/jw1FPHfFy
sXtaCRcMJNgSW0J4h06y+hrMqdX4LmkJi9bOLLKUj5t7kx889d6De6T+PqnIkyt4
ESenGEs0dDD+NOID/8aLm7vioRX8d7Q6NohcLJU6x5lv6A0EN+7+SJ/NzP4jFCNP
cDv0S2FB5/VmvlrC/dGWDMJOoZWzsw48XN4a5JTgNX/URaC0gcGbAB7IdU/anGEH
g1zvAVPSrISeO9XzfuQgSR9mZnklA+ICbQDLMRiw0y8hT5y0f5bpCPAplg893mL4
TwO9hlk7LT4lJnd6QByeYd0+jttaMTq9LmhcGZBJ8rgZpw+jWQA7mPE5BFeO6kHe
gZJInzOe6Bo3lP9ZEVt9G8Vpz2vlF5E7AiwzwxPsOcea6oIUoU1mkY/y3FH+P99I
anNpFtDYlNeFNkRll6Zkuh19y2I057Eg0BCN8PDbXxy9yQDKg6/YD52D8DpIg1CW
rFGfYhYikAg+6Ik39MZeiFfO4G10U+m3+dCWcVLupfoIXzj1FDJER6LDQh1TJPq6
gnPhaBQF8NxuFo8JH22a6OOOmIAPyrqmchdmELWV7wSZF6PdLahNpCTZXIg4TXBB
Xc5TUIKGxn5lZWFYe242gsxj5vp267oVmzy4Z5Nq4hUf+bE+mnrprCCxXXLHc+tB
eIDiv0Mx2InBBcnW5QjktlPuc4f0Y1cDrSz66KYwzmprzYsFKv4J2XrxFpTmJUCT
XHYj+xkyy2SFjmNdhCCSWabMuSSYWvYtXZr246hASrz3jY7iblri/bQeGBVwGqA3
c9rNnvvOOjot7M9ZY2HXJnOm+dridJ8Yzrn6/mTbJ29YBOywi7kJsXPm2WuOlWu9
GsFFmnMde5ZZhglq7862SIiiMxJb9qfjLPHAOur7w5aYqSc4Z9eP6/RGpE8SfJb0
GOVwxZ9QiXFyXr5RobrhZZOARQoRNTEdV9Oz21yD+Uq9rSYgMPSZsOx2FzFNeOeB
1nCWm9flqRQ6FeEEd6PpQF9H+VPmKBXWS+tDZE0wo8NzAIzKPNM+kJesCLfJ1qhO
cFPKHCnPovoyLnLpiGjdtP7zcO4Ghlr7/tQS9SZ+49W86zUiwBHsku+ltVrpQfPx
bB2SE4kyPXfvpiayHqIKsVBoIRDss3S2mkEHpLZd/pR+osdMD878kpHly1EUeXid
QIo26Rfo/4SNNqEntBvWAXZac98wwnlfqXPjgT6+EJ/QzEnrbbB9dgLyuxupy9s1
yX/XU6nsHritJ+PZtcF6JG0abQ8S3ssqtnNgIZYccpUHVOnjDnLv/slWEhZJyqH0
ZKyHDcc5vM6qhCWdG6n6v+bfCNCV6zWHIbxhdVzCI8Hlf7IgRPg4Y4GqKZ2O6GA9
QtKCJC5MVp1n7UjUirblX9eX2Bzs1ebmm/gYrM2yRAHFpuaCqIYUZQdOpmfopLyP
XjzZQWjkJSR6q9rZtWK4xc2I+KDG2tQSTZa3jLlUxUMk5LZKJD/JqokV/NLQvPd0
6JnJfX9N/8n3pta+pxTOEuWij173VGYNYgc81ZZr525qQiKNeXtfAOC2EvQ/6mnr
M7JAwNEhP31fzLRdC+ehPITmyHnpoTWLOCcXboWcjjrXS/eZjz4I5DTNBAmTy+Jb
F/7YA+EjiKHQaXs4+v6MdkaHyHGVDFkmbmuCeWv8/WmrlukqhYv5KAzjrVUn2MNf
EHghPwSzXc0shmJusakXv1Xmar7QUfHGmedNs06tLFCwFeB/9Ty7nxuC6g4DylXT
hKKalHtxRXQJtEpAfT+GSOr2LVg6cLHmink/ESYrMa1t0p/yriJ9PA/m2Io+4ZYD
Q9R/wl4qaWvqzGoULLlMk2tjhJhZapPBM22S4A5HNrNn3eoB3LhcSdTaTy0KaoIe
viJlSngKl+DWnJGbUP1CHTPOFVdz87SkfegxLbLN4v/AVXYYPaHR0jQKPmHJP0E3
fyQC+h/2geuypMoUx2tJay9/iIR/DUV7q3aVhNoUL91rdMxjVnDrfXECQbWCUVZo
vSidHMBcWJMRlm/IldmxwdRmHUu+NjHLpKlrTD3JuZI69IMvVUZhhfdAkqyIrLno
sj0JraaKZ9WvpB6AKuPnLG5kuyOiADY3/EyqTvWOGBsoolbV4J9ZZe+rCfs3YJY0
WljhGc5AqxttNpGGKim3gq3nDht+FayiLXrnj0DzTUoqixCBokbXQwRUm46nFAmb
jiQlBgTYtbINhtQfEzUBkiduMMxmHLtnGV6/9EQzDGXrRhtK1ZmtS9a4uxcDPwtT
A2xGZTQ+ch782IaomipZSKckGC4hYbMH+k5B5I1eq9j9XylkvD68f6cORpEu++NX
Yocd27/pvJ5mFu/F1Dnef10ldw6NFb7z1yR0kFVLoP+UcN169WR+EzmvKvpHiIGU
wU6ggdHDOenOu5bi4iywANb485RvbQox4AAa0P672Epi5cJclyjP2FxC7rrYiXy6
Wjk6YLT6LkuGvrHcqHuT+Ue2+gIenEzYxJcKpfhOlxWXCQ35HLZiAfuxr1FR4jcj
1vqowxasU1Oh49987SUAfTFg8iAZxBNWQfWOiEWlcEQdDcAT6JEVwP35uj1sEYE5
fLqICpgyCosTjL2wmnrhxcfZRzIAhMBsrzcb0TKorjEVTOHtQmeAkQ/yHXYXcG/7
HKgCR6C8kMclS68+iOQ+azuSxkgUz0KW6XtHelTn/emOCJp1w2QVlM+i+CP0eUWK
G3roaJBpTK2mjJ8oSQuCzTLoxMtwOCAR+TGKl7rkc9lvwEoM6DTmi2/eNYyXE9Df
g6rydDZ6xiFaJlDG+LiLd7oobT46YNS2WlpfC1pjGoxA11b4yMpByew3HUEkN6zZ
UCS4WYOXl+qgRWig+VEHCeVV9MbK6fohdb+o637SX3hq/oqOJRk80TuyrvGqLz89
7TUb8iGWQIFRXUZWHRar0l5WCibzanwyrRU79164Sv0Y1PoTlHfZRUult3/deZNL
Rj1kICiONjfyi6TLO3dvCFuXt+rsfYgquUlXSReWNplvzg/dF2iaIVBmsUUx9vRC
g0fzviLnkKoJ/CQWWco87+DkPKT1yq/DZjWhCDWAp1XUUC4FIa2hZB9MG1WXaCoD
NqfM3jaKWJNAiDEIQTMDJoKl/eKdWBZgwzlyi9En4qpW1ZQmYyJz/YqFKCPcmPdi
rDErLntwR2gEM0XPbldbJDkCzqzL6K7y3svRKl5/SCplFIBjUQ0q9l+8kLHNZ6i5
D2JnxKAATjZc9pq6q7MP+SfdutGq/+OurF1fZlnrpSvRsd9BRJjBMeVAStR8v9JN
jPTb+igjkUYf5ignpemJSk7MPfqj+NHP/7TyRacLhjkH+uJ4M1fNiyJpcWVojvb+
ZHZC+6nllN9ygHEomeW+x0rRQftKGutEykIm7Weamqe3is9PXGFP5V0lcGLizRzU
YUO8m/iVQCln8qRzwZQBQkDtaR9dCHjtNRydvfav+OpI7hL0sBAmPWcbQ32eHiOD
EUOTJj18eySU7su8RoCeKiv1Q5XtGDKZVY7Z7LBAs7whlaN3hozIfnWzB3NAe5b3
B+jSEjRMHOWSzPnk8IxoX3IOHXq6H1wbQcdHA1sJzqy3wAUFmd6ZD3m+hBQXhzFV
5nMkrF6dzCZvF7LccOv+ynJao2mDOFIWenBYDCDyt2C141KNtvBQHTIfzFl3QwbP
kK1rPBwJQh0LtrCwp3VU0Jk8xbLS+jT9onVxVvyv94a3VJMlnecrTCOzRRLF2hsS
fBa7QLn2TOVP2bXaq5dhT91pazCdH6AcI5/qKx7Dq89UragqUn8sGM22gVAtvU8f
HXpm+2vt85K/iRVCT7QzN3dz2HOpUVzimaX9YrUAlJdHiAgv1+Pi4UbijqWHXHRJ
8N978vHO32l74X3jqBMqsXQA84pgfj32uj6AyPH9W3q/2eLfVF48/APKmC27wBnj
PIopO+DZpp1oUrpfxZksM3kxu5jlhVHrf5aKsw9MNICqcx8IF+s5vwyb9J+ZAqym
9FrMlXZvaHJpVGgTVMaZW8DzwXiqulJpuQBOiydDkDq93+cs5vBTDJMXKlEuy3E7
aRDVJwsfOTztMKNTmvmNDdk/dov+cUf+e6aqaGb/v8X6W0pVkD0IlEin/7+/hnb/
c7P9KuDl73CuV7rENn4ZW4uJBf+6cMIERIMHTxPQ7ajvUtlr/KlsGj85RZbC4iSo
b72LNp1aujdouc9EwF+Na6ty/xxOWyeSfsb7xt7W7Xqbz5JtwYf1m5MeV2r47Jy0
6H2pMWlhNsBK/9HN9xOwKi8r8Znqte2lQoISuZlXtcjn4GJvhVFFI7/VepwXPB0P
lt1w5Hz1pET6jYW/xvlHK/b3mBpyJGwo9kIbVChPWm3wppaAOPVLhB4BFgywkrsR
J8RM5hQAse9FzBNdQ2nUmEwRxiCy67g3CTIzN93/4w7MhvviKxvmG3zHuvSwIU6U
OQ6glM/uryUqDeifu5qaOFboDAb7y5gMh8cEeq9HNrSma5UXfHcnLt5XjdX+NeMT
p3MEZvMII9dMEQZZUXdldF6xeADG9JvJEVxUnUDpAQ4mZ/BM1Mmh0a3sQy00tdbr
7RvuHl+zqc9K2aAl++zhRMa5mNRhViD0/QTHPH/jUAIzVl4hulub8qIkZaFEyG61
QqfeA+qLe1nOI3I3hrSTsun4WIz0DJFc265QmKXk4yf5zCOlad5OsNdtikRY3uys
LQyLOCLar6nKf0G0U/6vE+zKKsM1Nyc4yKlH+PUAO/eAfG0nKNaQyo4PcThxeYJ/
6y9Z6975czPqSZiRGKWRAGLdeGyJMi0qx/AsPb49l3igk/gWaWEyZQxLU4iiSNRj
KlGXMPMgTLuMlDQ6FZPkXl/RWRTd2bdxf9fDikLdUi78uWFt/1Zb2caqZ5iC7hlf
ognbTnYUpnN92YmkbTdJWIrlpTU4hlgN/N10kx5QSQebb/jx6tFG7nT3hEoES2Q1
7u68mDiD5BiG2wuW1J+vwBHbC/jMCWrL2IrK6LrXAPxNn1hcYL08Pruo6zZBEyS7
V2UTxX/zsvAtg80buMoh+llrFfJcUlMBVbk37Ms7UYLN/iscn97SrDVhZj46M5yW
qsABLgvJdqIHd3cYcIUItJLNkP/PZ8kyulQ7TdhSHtto4nP0EeGb6yHls+/eOxun
0Nyun1u80rK87n58dsYV/aq3fF98pMZdNENwyDl8PHqxot/IUey1XyWwtYoZ1QqS
L/spxohcrje6XuqWW0U4regr5T6fR7HNyDI/J/WKiesu4D6Ge2VDARM/sQN1cpSQ
GB0pew256fHNB9ze32/tIvPfYSUzOk98peH2PV0ey0hHrbdn9dJ+y+3yciFeSzw4
UGWyC3lt/Me2uvX5EivBNfgkhMCOq1WnoSj5He0oHPwJREWZgmBPkEGw28b1Y2UU
KVeY2bVVxZlreDZU1+OKf1UUwgb/Jt4WaoOJuugQFjteb37NG5aZ+AHsNVtXlS41
lSiZ9fHu9Xb15jeFRQdzulHdQeCnx21D5SttT1o94WE/zBonHQGl2ejjLZEbUzH2
bEiKWPrJ7p+KxKxwNaXiWea3tG17Jm0Zud28IB5hswIISVqQxAEnDdBdv5V/1T2n
xSR4o9QbDzbhHUh4UWZ2iPs2Zxh8uYbVDtNP4STAi2fxEMtOP3ulNDIyOevIckIq
SL7FugEz6iPrFEtQNfmuEZC/A6WKuHPyvKuLdO7lvgvkrHEL/FqfzhqLp5Hn5aqW
HeYQd/pJI/zBEIUqVR+GbVjkzxR0IP9PNxvFGtx8YAx+XXs8NuuVRjd4WM8tLcwn
GTnXzChF3TTlxcw5UdyMxHw6cmc24LhbvZUTC1QWy6qp5AAnKjEIqIPCYG+OJuPQ
K908Q9i/luP+aMO/yXGXTtOipryPAaJkjaa+VP9LgUdlTe6lvI8WOwRG7csGcAPJ
6v2VLM0+2+ZLo/u6EtvJyANqiDmda2XFANQFJgA3rcLmw1UriTlJqsARUZ1Z3/bg
SLQiMOrWQBEGVmOLot+UsyL+B849ZeKm5ja+Q9OHqk1NUhhVBQT/FjwmWsTjYYlS
RNSGRlpBO1WMkWke/m5CBZTsYwOFdq9JffSUJBmXvhN5b+reNJnSGn3m9S6J89B6
VxilicfcLuupGrdLOVS0yjOwKqVekyqWzyQ2M4TFDoDXcrSaaB2HO9B0ZlvjyCC7
1/DGGJYzHOPHgyDDhPHBMHUj7mr+k9Xh44BQNTY/AvlaUDC5HjzfxWMjKZeP9DVW
DcwXAnIPp96wpfiC7i+aqXmTBMW6oj/5YH2A83xUfIT4jf3gAB8rySAld46+EVGR
oddE3SZDsykgahdW54r2TyZLer+u60rr1GEONITmkAYVbHzY2GKqRajsxpcTwEAY
+x0SOXPCDyPINs4XOb29uWO0GpAgsAMALErJabOa5lmtqCdE61inNIGCA5Updx0S
34sNVSbzJ1bdTtp+0ZSfARpC1LDdZ/UcxAZAWQOwYuS+4nOucxpTwCW6JGvhYQQb
3RIomYR9jkN3ZwFUi/hy2vspRMF6zbUxYPBawWddoRzhRuDdNY/95gpOTi5hQw4T
2jK4gvgpr3/K5SAXSqJcKiT8czTCvtHBEkPDbBSKXQ4GHFJmIK8HlA2Knwe6SlU+
EF7Y0gOguLO+SNhokOIsjqtLBrjPSFRTBOZ2XbkyuuuzxWpHE4FsjoJ8DSnuxz0f
lFrpNSPEhIPhAEH29Z2cBZhma11FYP2arHvsXLs4LEHhBba0SQw7YeSCETxgi/mI
803S87z6m12h1shP6tK0SIaC7LzCFy/M6uK/A3Kehx/prN0ATeLYgdxSAPWNG+v8
p7H/JBp1Ui6Lw8a7hOK97wubT8gI2d9T0InmWmvjEzk2olc07mMVuXVn5+5d5bRY
XMnyughU1TG1sAw73XZXSE9ZtqfsjY6AuUFqg7ESElqOyOvz9A/hMReeA1g4Pzz0
jTSRmHK9tzL5CoZZOJOXFQp+wUifxF39jCHShF15gvWKAMxoCpBJhYhap0HeT3WL
iT0nvN8rqhyG5PGmVS6+Ws9It0dGhNUrpemq24ZLd9pKjyKSsTzJlAUkUv/522Ou
fIO9MQKL8BqS/4TUfGSDManCD6qQ+BIYb2XB997SphzbUaAZQWcZMsZITSyzwWAS
4zz5Ai9dhzVUfU7YDgjV4xvYuZUZQyYQ7SgvzD4ozbW1/XdOA+AUKqCMs5KfM9y9
dIPZ32c2YTW3SSwLmiWqQws5/uAtwoGMUpmcXKrCEoJHR5DbmLoyakzsSBxiPizl
Fai++VxjOMUqvQtQzeAkuXMAWIdSuvTKvM0wecRobyKcOkUX5Fi+QIXHZYKN/e18
Ym3fJuF0RZIqZ3I04aIiwrY3AHrVZ+X4v3b+pXj9oP7j1UOX6avOpf9lE6ASe5Uc
Xycup7k2Sgqkwp0qyAmCTFWn7bJ02pTUo6VDZ4LRqh0ThYjIfDeL2Tg60u2IGG9T
BpsR6aIsoBJ3QzlpgPwkCPgP4VN5K2EKyCXZr1tgYf1GWUIgNE3ahT2W2H8DGGnM
UEGuib1o/rIElJ2XleGtHXnWlSiHUz/N4ekypHZazMgWEriYtyVxepDBDodoszXX
Q/vSFxH8Mxcyy0Gb941QX/xro6fV8lVUqML7InVcl3U4RagTlI8zjB99Gxsl95P0
Ia5Q1PDPrkZYBbrrjYtZpKM26IqvFQ3OxLuEcjQfGJRESUy/yb2gLqIrjZWAIS6Q
Q04Hh14m4/HEnwUAhXx8WNnkFO4uGccB8QkI/biOmVT6k4Drd0uenhCjDWjKaA8Q
5dlILbqhjlLXujZ2EUtlBx97Ow+O6EkeVYYyN76Xlkbbx+qcSe7VPMRrK6ZQd7bX
X7iOu0Rr8IcLqdxfoSgf12/29Ivb5EODSPJL8oFaQXdcsH24EXV6j8CE9WbRIP8x
H/HcAGk/F9gpCjfiutU0NESxrqNj6nS92mpm3SYsEHdhscCyk9vTzzPCrfnjTWn/
Aqmhbgey7g1/2EH2TVBgHHaZDHtN5Almj+8tzITIKt9IkHT9Cx5ZbtJR1Kiz0whL
zEy+qw9FfDVplzdrxK7sqiw6qOU+dZ+9R8SiOo+XMyxMYaNM1qSPoMH6FBxNsXAf
Jubn726YfBSEZlGORgfy3z8GBif4hA1ZSDG4ERYO9RUFoIWQxP+TS8P0sJ9TwqfL
blCQklIDQN1cZYgZiR+Jco9muiOC7CIVZqG2JmlomxBBgM21vdvm3LGr7cq0DT9y
Cn+D1LHK/eggpOLxrOjaoo2y57/yxUtoiAxqEka4FFrnqZSL397akquB867i9V72
65/IRUrncb+CnE0Ztfcv2UCMLuY7jbtIPbsvKOoXCuNrwb2Mc+ITamFb4OhkGIiM
VZtKUmR+WARZ21YwUx2D6nVULCSfWIpgmpLEPeGOdKjJhs4Lb5uDlthLniEvsz/P
OLsyNk2tf+TanSnT+drKozUPLIWudAlYcYamFE6Wwm4hY3/7ti9NuFEQCIZqnRpb
LTpN4+KsAj1dd8zcMMJmi++KwTBmLkI0KjFQGzqYl4ha++N5kyxT1r3lB971yIS+
6c66a4EhbGpQLtOgyQYrv/pRZoLf+lcITv67CrNOBe5QYlYrNZExJNOsJjPi5twP
bT8MniUNj1zAbcoMAdysAvP1iUIFYL2RKwEuhXvW8/3eLLWiiq1DnyyKMAck9yL6
MXpU4AoDRJiljwGDLv8VYbff/KL1FyaK0LgRShDe6zt0qW12RvnaQwUbZHdUDPSB
Lxh6cMdZKmX8xgoT7qx/HTE74XTM501C5F7K6Ia71MYzqfT1vSO93ucCMcie319Y
RCfhPbN1iRN0aogu1DhX2YOWvRFOXuv5GVIN0QweMRi5KSfKlTDpqtZHJgNkoOYk
4Sig5VTKdpl0Rvu1uVE9bRzjFv53CIbg6lGw7W4UoZkQz1A27+20k1JB7SNzaRLQ
M1HBfAiRw6dtncPdw0Gh5YrdC5XlvHlSDJojLNM9yna/lYtG+Uaa/TcxUFI9e9yx
uKquS0l0SupQaoi6Pn/ynhuFwQixEH411U9XymJPlOu/Gr70uQSn1MnQNUGgHF6s
4UqVCjPudY2CinQA05bsof3Bq83m+8E9NL4VSsD/7SN/rvsJzG2+aGA7RNqnBDTM
qMrqCv17pApLum8ro2jLekb2G7s1njl/sIvaZePZpGcKUx2xB4Agf6oul3gCMbJh
LZhUhFGWgZacgIIMnYGIVktrhPYfC8g5HHeDkox5kOsOkT0N21O3nBZUYqGZpPiY
FBMlYh/n/W6Xx3WEaOeFV6Ss+mt4VWK7EiJM9iqehvtzjjeYkSXeuM8ewvnytjdR
m16k4nppzhsk2362uemA/QIGjEn6hXlw/GIY6rppYnKHS6t/Q2Yyu7L9Nev5C4ak
LX3ZLUFcOLZFvUytMGB1cCl5CU4MIFCHkNLFRbDs8QiinG35HmfdbHRfMeM9Bn0K
Lik953MwZ1ofBtj2tqob4wMe9z1RDL3R6LwDUJTkaA1RdiOkHzByVgtwwcLviWCz
nVpxQDl1pXmk2Un9NEfRRb206eUffPfuOQaDRQ0WID4VsFYVDjyUsUEBnaGO+VsZ
uE24bhDRT3/dAdhO7ZViPlh4DDWuXa8i6RzecHi7k4B0G+jvltvVDHjwss1g+jHy
duPiBL6lTuPpkNj5EnOzlp5lT5K0FgOGFTGSVxE+ySRjMbwD/VB9w72TbHMUfcy6
WWocS1gJXl16ad8pikjkd+HL1tIbQchobdi/f2H/I9OoEo6Y4E6IZ0IxxN3Q5gOD
9qhM3qPPXjOrqrbj+HzF0jTGOSpXSabYpJCwaLZMs/pSAEXu5Fn6zwxX7pxnYmFB
BvWb2K3DVhqYUL2qeSlk2jsaQSLzJar67Ht1by5EfhuT9yMh6B/GDFLe5DTciNbI
ncSSvYh8W+bAR4NHHUtODZT0QghYpgU0l2usJrvuN57Ap8lkyn6hLvECj/FkzLwE
A1N9EmcJg4F1CrkmC+Hp9pPd394VAq27LFzJyPA3E7WAb6ivvHoXF5xQ8EEUSE4m
MgFc8Cvp7UG4Pdpd5toqfrx2mZ5Evt/Qy68peqLm8BuZ5pIJYwPGEqlYSenOW4Sr
OqmtyDw1VI5bKPe0Cn8U+15BYpb2rbjV2H4xNq2uydWjL8efmFxWyRlT72ztEDZx
kUNueTOazVd43yOuWQeytClYObqAMOv6WBtl22K/ZZAt3RKrMWFWOl1iQn+Qm3d/
qxE+QCEQ0fK19NI3i/0iGvQiDMS1BbQ1BjMxnE9CU8Pzl2wpt6xPww1HF0HEC5o8
Ok2/1zJ6XsJU5UO7glVOIfIgUiuz+9ljPujTbOC7sQQjr/9aMSWOT/mGgyxzua8L
cxs7FPhN28+vnMNSj/5ktRLKhkMucOGWJLX9hcDwMt7XTjJm/ygMMFATBl/mG22f
mYchmAeBfIBTkcf3kygdlxf5twWtJUsu+W81rVCwS8sp01ev/9zBeT4+twz6nJnm
/XLWte+AZk70OqsYSbTn6rWGJrTEoIPnli5HqfE8vev8Pti3IGQU7ZkrB1NJ8GDv
aYTzYPyKF3PpT6kXOxBvXXIcto14aqT45IQhdW27DQlhWP1hsfiDTq+zG61Ra1QS
9rZsd0fc+qmFaA/KxW8+K7yzKocDGy/SGhOOqX1nOEWIe1sVQwR0Cx7paOSs42HI
RDfUrYtEDHX/CJyOqQbFd4E5TKxcSpcmRNY3tUn0RYr0L2uwk9Y9mtMvEyKdWc3Q
KzYyUwPBktRa49w2kllaH5RKxTGIDUMbo2+OBiL0mhLSGJNW1QtgLpqgEP6OUZTy
O5u+RlJFko5Q2C18TiX+xPRT8BZ/kF6T0W0WQ7mYaMoi8MH5xRvu86CISNPyzjFC
iKMoNcVYVA6WpbSJzJtMW3UdLIIgSt58ia6TL0/cw+yUFPyqMwWbVg22ufHLSbYO
KIe/ixywqj70eN4Bf84/TEhKBTFZYY4Tn0+YlSqK01hFKklI81xTbHylZVPR1hYE
1pNta1g7mfQkJIYdkWNwoQPC24sK2Oeu2dkbGNoYHC+lWchBQkFGO2W951Oc8PGJ
sqtw9yCYKk3M+bWvZvaDrL85Dej1g1DAgO9+GCMutIpyi6uczCb2KPyI29Fp5v30
JoVx3HbKLxHNpLKA/IvSxh3Esgs5pdzZMiqCCpmLkloqD7ahbMCVkr1qMmKzsJMy
vhGD2ezfIshCTybcLH/LR/PNmPtvBAq918kUM1QS5+f7mjGk2js5SkOiQAEkG7fw
W7OuwD7rOpKNxXaBzsB/zEKnMWY6Pf5JKcNjhCvsF0jo6Dz1bPSZlMKVQ95n20af
98u24Wt92JPmBYKASmPGlSUbZwj9428oZ6L3LkQCrHFuhi5sK1Y+Qnc0rPLgZWpC
U1utA40Gftg0GlViYtWYy8tnySVTO3SYd8q3PlWjgWEAKJD1VHgqAEO5BxfvnFny
6hA9RZiNtrh6P/VaDICZAqbK2zjvHZcpYkens3zgOnEAjpBE5REeMnvwQUQCbCUb
evaX0wovFdxVfBjWvVGfD2eraDu/ftM9hj4PlEzPGOj12aSscvRQSSmhjidU20Bd
0+IXzReWYkvmUcMmsXxI7Jusa+P7lsJ8ldTMKL6UcRJ9Al3F12NglwArDexunXdt
jaonXg25wNhOqTV+ju7PrqRLEFPh4jL9FrRrgjqROoZHhZ+eHljva4cSDbyJwEzv
sMtKYhclCubZ3Yvm5rPTJxjwlzdLaql342IlGAFMJdg9OJDeBCS1SG8Fawypk0AS
MHRLgRii3qOqsmMaoi5l6G0oWXnPySE0/X178t4tgzuZmYCGjVYXOWF1FSPKygR1
mSZZiw8lE9hd1HQRbVWBrwhbPSiKUTgj//EfrCySiyfees7oCuEXGvpnl155OTiR
uXTrMeprg7cr1E+/U/EyX0kdxsNxViJ7NJcGV4A563N6JGuvwZsgsV63eSETr8Zj
UpMSDWGQZVRpizp2IMilAv8ADi0Zj7C8bs40+goWQ0IpBvZgKG1iVfpjqrfVZSU4
I6fUVWJ/G7okxv+eSpBeWN93H4yDAxN2Y5jM/B8mxTPYskXeCaRUjzFaGnH84SlZ
i8TdtHm13LfV/R/9sCuRBoWtdrwoLQyqaSm+SRhI04sRMq8QtwMztxNqnje0Xi+r
ZKrXbMrCwSNeYinNy5Mv7cfBUSCv0dJH/kHpnfoA3/OtPM8mcUbvAGNR6+iLVGom
3rDpDkA54liE75PHwQDH3AyUgf/KjOda9Aw6hXSTKCv40V++4UECWFpNbKVzUNLS
uDln2zpudoLrwk9JrtBdCOiF0sO1w/duK6E+sbUL/0O53K8lvXBzTUwS6zPArkLt
ThL0KR3Y+EMdH8OuK327TdgrPfIvp923u1pGkc48toX8ED2Mm7Q4m0/MvACcCNqX
fWnj4c3TxeSlMg4LeCwGpYo1l2rZY3IesXfw6gCD5V46j+yrj7LIfoQnyt5NboJm
a26/htHf7sekDaRXk3TUsYq+K664UxwpFxzdGL330emvtg3rtXNcaKaUBtK6FiBE
cEFlTR/wFUWQLSEuEKnIBFj49Yr9Ue97SSW+LIajSTk784Myl98Y/O164Vmfrz8y
PC7ZloWpDMykp/fAn6zPcXMIXg2zeKtU6v84ipXZQ8LkTuLq32EWuhOs7NLOZOPV
gFpnXiP/iq+n5OKm4osEniBlfVr3+4zAdTQasWfaQUQu7JLcYFJ7e7cuxzyPm2m5
QFpRFb3xEGSIrXCbMmi4CAW/oSC85cXvxgNwEOPVMgMwFizWvfpPQdaEtO5yanct
lvaIyoRtAaU4EcBHmvGWNv3moBO8b+ekLEx9VSfTANhvj93mabhqoaimmosRwubE
hE+rf5X5+QOUj3GBOGVpzeDW2USS7mnajDg2ccZxDyNOS8KrrORzZFoI62/4bM3g
83XTElHwaf33Q8XLI6pKswkqdUqNQxw6Kpv1Nxu9huxuR09Xy6yKzcPp6LSunl/2
LB8YNX7xn+fvSS7dCM7e0Jhalkxbm1VBG9KWjyxrEk1IkYiYqeVFwKNlyHM1bFgc
Atk2RtoGbrt4wFpXCZTjV0czBoaLjaQUNrWJNHfQKiB2MARHEzQfECr+0PFqQIs0
fkMuuL6c3ZzmSE+wWzGF5U5AyK6T3JD//agWvkxSz4y8TCEYEg7uk9Mo8xh/tEsw
h+rWL4Oyg0mOIjLcltpDIovYzQwHoS3N2WEbUGg3laslwX4ZSY7VDHfsgO3zA89g
iCSgRIaKOiGPjWB8ewejOhpvUgBg7YBJ7lBI3lbCltkJ+cmsWSRX3NkoPjf/jXKc
N1idpKmnHoy/8DWbR1CvQGXI6cbjIC8/Uu8QbszbUFUUeO14bVBu9XksmvQ1IOxH
+7EFBLEzstCN33gxKA+0ybU9FSneUKIZZe42gxa/EYVPOLR9AZgGzBVyZjx0tzaE
jV8nYaItF5XCEFuwH5IWwWYLH1auIPYKhXNIvWF6tw2qYf6mDXMYB0KDPcwMJmth
Vzvz+PdqHzcrga/jT7RSO6Nv+gymTS3pa3y+LLfUiZVXn7EFcqH3+lLj1aDDpNW4
Rlu34y/+lXgnIG8kNALc0Z6sap6KHn5B91nLIWxnkhTthA/W5Y6HMqHEmJPddH3K
U69yP4DsWKz2T97PODxRdk805Y2G3/Izz+LTcW1kNIAFLfGQH9GZABJxBsyGoHKC
Zbhsefgv9qpCUC+slbVYDGEWzoLcrpl67ZynTZWJVzKU9Fu7KtbH2/kFt7SLrttU
vOEO58HTRaqj9pxNT60vlt7HOcmDKSXGn8BVPcRnzR9t8wjdoIk9w3Z3h4bWbmkr
XOelq5nh1v/qcb56PFSGn+EJQLOKtoTfUItzrXeueoYCcBvCKoIXFIAzra9aGGlJ
Gnh95a+RFdmrFqL6tewgUQZxL22xvQoK97BYANa6bORXezYYcy+jLOBDwZg1Vo5l
lcj7MZ+DwXHZjezqgD8SE10Pk4xZj+KVbVohoiPbxEi8tPUmzZ302uMv3XfV1Rhl
Bln1QVdDBagTjcF98VTmK0byQXREqzVzD95iZOH1EcqFfM/KnR4XaDwwnGaPPdYE
818F/zWYFecPI28w3tgDg5xqM1yqeQPg+vMms77iyosi/MYTw8EYLvY2bdT94RZ1
trajwSB+prK++a0AF4R5DzGW5tqYOXWUVRcSOCgI+5Gk6vMme/gNVclcMcXBt6jK
Veizy31potl7tEKN1iJU/P2lmih+4izMZULu5Zem+i6bdvfvEEEJW2mQRJEHUgh5
oVL1XT3pP9GOBtKdjgDuKrxLUSWbOnGBsAnqM1l6ysunTEjgY13FP1bjwcy4Blb9
hx4Di6iPiI3oAKHNuJQUsjpQT/6SAdJehBGOq29RnS+LueceajSXa1GcEXDXlMOc
agiTDqRfbGhXlx84jahewWcwgEiyo54EbiGhaVpNGW+gD9p9plCifSnFdaUdcTp4
bGwiEjHWTqySFMmf5TEc0VxRCp8d4CT3mMUFYO/Z0eNnH0CX5yQn4uzF2nv0C4MV
NS8CzlDYOPIxuiWefvw2t0IwT1VM9PXdJ8NZBWTZ3UCpoM6LxQDNQkj2j350jhpZ
OuiO7STZx+IGdreNytzczVSQrI8y02OYAZ7yctCzEK08LHKlLZp0Jd3MXJFUnETX
cuIPtrVY6bSUojN/3p+EjT1pW9GDIcrP8k/MHfGDPB0Oa0Whu8O5llmdgc8CIMCg
hkyygja+Ao9HrD8+1hzHiiCYx4HLZNzUTHSI9uQ2cVebmmiHIpnx3eySb/wKVjVN
g789QS/bot5JmtJey2Lhe5TGsmGsM5tnDAfOqHEdP+YqMr/NR68e7iOZHfd37V/x
biFYpFWt5OJTvtoLo/S72AxEFd9MVfdrYtcT+tV3x/EaRUjP5tRvAe2WsAa1O2fH
1xapDaXqPsjNuA7AMH4bvKsyfsWV+nQNXZ11saDVzISCpVZ+EnGoZ7lJRTzaXh1E
VbgB72+XcZogH3dPV6mY45IQRtW7HzrNRl+3KKps1JpFVyXt09sDup/VG7GkmgMr
Zi9dSr7b5ZaWNToIZwyDBn3IWpU1g9Uyxn+9OBmxdF+IXUbVNHMYb+R8H0ZBH0ae
3FFxci3GUhL+OSjerchg5hp0e26uCCuDQup03CdlCjd01UxdqNnneVY4tPShU6a0
ytpGM09+Ja/2Ey7xvmSCp+GvHdkOrrWKdHs3zZLO0vh+ld/DXd4eXjzJ2QVHofZy
N+Tr5442LU3hj84sd65HXOMLDErMEP5og6TZtRzibYuPNK5VURzCqcONfBh+uSl1
mly3N3bftOMEHNfNbyctgUCLsv5LkPJRUDVRu7oojkEeMmpFk9yHsvXj7OOu06fc
3hMF+M7QJf4HlKghTEuXOLjON9YOGa5G4wJfb5HNJ57BoTKVlfpYMW0oCw4pi6en
EHsR5fwWhiEMpD+EUTuu47BURTPJx+dH/fcrjfmOWDxz5N3lJXEYUfmeuK78klZU
F9TymFF9xrrEZPyDgad0eZebiWp4/19rJZKyqWh1WHy419CA/6Kw6nq6EgtHnVcp
+3vZjPJ3JhXoVLtF/jV7YfZLj9e6IvumBehM6bXCjZ7bBROnGAPuURXcBxStnoxY
QxEQGcSgWPZnNpTqtLwkPpCPNPKJNo/J+0Abal794pOKZWjoZFo673LTR5/DYROC
j4eQBKMfFYw3JkyarIRXHtVI8eMj6I3uOxCUXk0cDGM9N6oJQp4lmU9cYYLMZfM4
26btxbrH+tPG7v1xNoAfdXNLmQvUHl7uit+Yrmu1zbJfjvrLv2gNXXyNmZLblOxk
mop/bdgcWIwdVeCCkhi1lt+Im2MRusgH9+ZkHhPsTcmvG/bS6D58THdCooDUjKbK
5wLFdybinFGMQvzP9WBng/xnt9RkUBcgE/OJD8nz5Hoo39iKjZEiTPvFB5oPR94F
UjopCZpdzQifLdsO6f7h4HFIVNKuYiX2XMqTIPKQyaHt+McslQ0MHFpNtEzLWsci
VNaOycIxzeQ8opxM5Dknrhl1NQYGM1oi8+MTdnG0ACXx5y8TYrPPOHS5rbnWu75h
yML7PhoMr4sT7JIPCUEzdfchzI5Hh/nmMJ2Na1myWtvp1+3l+IvC1M39eyaUnvDA
nnOZnXmApDpFkAjNQwMW5hKGwVwI7p7+AeL3L1AdwBt1RXgehq5hpdXoJP5u8l+7
DcBEf4SAy1YvlAv5CSHZ095CRBFOFTb6mno0rcNdWMYIj/6AulbV6Eza5DuWiTtl
EYdkMkYhTVi+V4Q6lbb0BohyWQZsYxaomcg4Q47cE8rvq2LDHIoG95HzlK+YY9MH
nQ3UaHsCQ6x/4q+NdjdMkDZDXa4hbHg73DAH13BX0SHiOVLdbiKv5XfR+XogEk4C
5/2oxz5oNJrW185BE3oYTb3yoTW/K3/OyksmDhF65OYcCUgmhmnmuXgURqxHHhMy
ay8zbMPOK97SBwygTbVoxq6chmh8iqzIkic+PB2LOHIN05BK7ouB6pLcsyi5M+fo
mX5q6pW+9kA9l7+7O09Cafrs4qOhkFYAUJcCxyPJRfKmjZhdrwSXdzzg/iczo/4D
/bXVqoOMxEQxPcHVzowgcuwOhLFw8tctAIHXhEGHSHpBiBxMiTU5q25Xx1raKopP
QhZacdh3qPiSkBFHsA66Oel6cMwv6JFCBaQ1fTwbP9KikMq/SFdUL3F5lBDljR04
VMWfnMUi9iSPym7qmKXUcGxfuRfpCotAz8LHMz9pQ9vA2eKolrQCNLIxwMDCVfX9
sva/L6+qYg37RClTX0tFGe6CFNC1O0iDD4AoxeFGUJhO7sa6HZH7zZKvnPDOWLQB
2+/TfPwR9NjsSEXF3rlqXSpeVlwTpB05U5kfVzITlce9r2+J4qAvlY7MI6cCDb3H
7ISpS2JihQgm5zb+zKZGfnNsFE0Nko3xwUj/m3QAn5uHi5SC0UV1s6Vdhb1wZ0sp
Us134O4ZkPGKMcyUD6QpER+POCYJDpTF1ZTMM2O0TklUU48VfNQm6Lx0fX0zFi1H
XffIGdFfrb4aq9fa9gwDC8D7Mut1pjbIpfZ/nbu0goNmsqGqohTQUtHjLClsGb7D
acQAqR7W2mDJ4klIkBlq1N7qlzjMW1yubWP88fzI/rvrBqygqT+GJ6X7Kg41STzF
xMg4EqRrBcxIiRfW/CFSCqnmwhZwH52Jg+vWKMdmcOJ3raDiSu2AnoDNXRbSFTBD
eHru/tuhzZCHoeuXeR3gEVVI9lFnjYstbnamOnWRgTNadmvI4navWp0EFg4pDEMm
q0UmvRop8ybxXvaAYinI35UTE3sg7++pB0QIo+U/YauDASQbYqD8YVw+hLCR62U4
a2nw++2cOB4q4C8/2V0MjtHoTPJIhej3Bae6ssmsQb0XSVcdVeaJUBvBb2/t7k8e
B8M2hHJbIgZTviNNWFkFoD+4gChAW8/3lpjG82luYIbqDkgeTJz8XiBSrt6unXCS
Vyo0vZHsrXk+BxE0GZO6glENM02BMBAvn1fT3HeqYde2MfuYhXvDJVbfNVj3yGrL
3Nz+g/PC8FMstLT+tzr9XrqWUCLjFY1US1tvHstok0uV+RuzBRZGk2EQu0vc80la
X82CniMA5OU4rm5jqlhsYlGc1jAdNxmCYPEoEi7cS67WN7Bw8oJVY7XpeptwMp5f
QFWaWC0IaRVBhmpsD4Y0vtvT91YpWISYhh2IZDXQMOlLNOarD/xkH1/CI16ngric
f2u9sLCeNSjfBBsaWZWELyS9R+r7norC/cW2heuUDmOJVwm5tKsNlQzY3sYpNUru
IpmkeuMN7tCyMci3+rQM/55B5JAmalJtwfLHiJ8qCxdn0fnRB3Di3Ps/I3kx8Obo
D+ATf3cRGpUb4ZaqzlmhG3ZTAr4TnS66/92+atF8Qoz209nJ5LhiLxSFXjY6VW3f
o6Oxk59dnI8QTraiSwW+c/FEaUTC9FmCM2VlEDdPdFhk5u2OURrc4g2Km60J3/FR
jtgjuPOjk7v65Jv+FZSwnrPv3hVFzBa81dfKTKAHzeuX/rHPOcJGBbRoMRmYHU0M
IU1tXZwHwhxXr6Dv4KYWurgm3V5nnEcFlTpmnkGW3MhdqP/eL7nBhdTEZ8CJmL5T
Sm1Ly2K7JIQgVuTVJIkCLIVHCHTUW12hy6pG2MPolMQQP8KASEuWr72HkCYtAZYZ
abaU1z0ERjgWJaYsRD/+vWGfWDCBJHIc88mH+pOZdfU1DylS3V4hP45JYyfPq979
VN4Tnf5Z/aWOEe2+BSqQNMGVozuDN13gtyzkaDznxKte+BsA3s9oyEHy6TpWH5pI
1lHctAUtWEM9YfujUyBd/mGXq2OcLL/cnFD/doL4Z0LO0VOD6heIrCOyzoI+V5CO
VmFHMnp87ilQRaSTOeQ2Y9fJyLZByr5VzNCqHiS0GRieB9HRvadI6G+fHGp+Rinv
rYps66iVPAZ908p8O9YdOMtqiC/I8N3YgJGu2sfBzK+cRTaJWGYXC1BdWxclzoYk
pR4GHw88wxnB4vZKUJxzdTte86APP/E64igFZerNnB3kEY+uhiI6ORXpwXakoAPE
vvVF9aQLkQ0yZaGX6qSArgM2rYmvvptu5/Y+q0BX9Ap2eC+NpjRJraUKMMN6JPa6
zU8g2fC9u0Jmbm0+tDqhtVJEU77zJIUyhOkOb0vEIuS0pbbgGK3lkv5dMaiD3s1T
NDR1VHuxQ75SsapLCWFF1EAtdlWy9QTQ8GBbKs5ir0Si/a9Uls6xy/gPpLcK9jNy
37oB9+6YSRDkGL5ZbvQj9JF7zYLEAc3Z6HCWkQBEjVIaPcHi/UEJIjrGxGN3lRLU
yRGdlu8wkKO3h9idxIJrandwKbCVhs9fLxsq3URpF0EmP8JHVruVGyG3oj9fJper
qCfRs11MPrfUIFFSDthdy6Wy8vK1SB7UNMBY3DzaRRUnybImCWDlPsOCCdJKP61R
+eIkFMeTNK1IYoMJ3dSoDFRCFkh1q5JDRo8/ep7Hl55Qlu8CqLLLF90GOlolFNso
2h8zZAI4nJf9+0xFZ3bVZ1toq3uUq3RJ4met/e/RlnCvRDh6LgH27RUBLpMzD06g
RYbcccY417YjO5R8Wp2MjD7Vtgj1EGzLoSz0Nzw2J/NSEvPFruz1zxKAyT0sJNwy
RXGQ+3BhFtH+SHDa+MNcU3WGqM7RYBg6M0Ic0WKYVXM6/JbESmH213P7ckwSqHYb
77mDTLLKIRW8mkWPVYK6Lw/1qwYCxB/jumwTn9qOAtsBQQFfjazhcaR58ANVDzTK
f7k0rdquApxQkdeAwROMY6FkVzh/VqMspQzeaNvMeRwZpV5Ag8bfVKeTqWYQHOCK
PemTo/rbD9He9fwIMLCrlTI6HZbEaltgQCAD9l+zC6d7QE/TYZcMbBLJD/nzbVGh
c4PJDeze1zc6/0RNJFgfYbVL3hh1oqbEHaW7WuOkwLkCx7SuPHYDXwUGF3e9pAKH
AC7sE0GLRKEcPI6rPAuza7CVlaOfaY2iYstdLwy0TasfYQnp4xnln3zAB9Nu/9eB
fPiqLiGrTk5UL6tSzTnV8aevz7XlWzVGhpOhyn8lLnzc1iI0sDJgTjRBIByOBiW4
JOjpRKJci0Y7IZ88Z0uvlYTx0OJxFKBXdOckmRMESbISA+px5SIvetIhymfVvJSq
iBKreorpINSBp1d0jlAAuKRjhYGUWRj/k25jjrp6Lyb9eQqcQWbPPyHvnWPrxR/w
+Lztf2mtQjb9IIuVKxJ1TffMJkyqJ8AtEzmShRyLk7NtCq0t/OK6pQ+qC0swInIt
9NDM99FlDKQqL8CCkK46bp18tDyyptRKozPFuEon5KF16GxabgwwJ82y6+kH8g/r
a0t4E4m/vv1Tklb6zy4l3fc0VTYzLveuvxcnXOtXiI8jklpWir20wMIvE9anykLk
loamKp7Ws/XYANqMbXSFUilpFhX3ux1c3pVIlpxseqdcA4PV/7ifiipJkprZGbD3
c+ysx+X1X6XWx5CuJfTBGCoFiQUBVwOMwizjAiq3SrDqZDpkKZcfCR1hNXWDx/vd
oexPTV3imL7RWbLkf8U1Ijkn3jXNEQKed3LI4QbGwbflEAk2iTzeyGpQPwHp//2G
zbVfphEeZcxe9MbfI9WxeL6visquj8lJRFmTIWmTS7gI3dSDJGvv/Zu5ciKZ9Sjo
61QyFH3lR3qhDjD0JtnqL4wLBJc0Y2JR6T4q63hA5QrKiaPBWYExUh/ZD+QCCB30
OZvFbj9feZDDKx3M4y28QrOnb5NStN+Oem3ZlgkVuI1nfF6cL0q5lyM1Vg0WcsZ8
h8gfeN67HizbmcZCyfvVp3+aF3oJsz00VzYdXGkc3ZhyAYoTH3aWZZzJzwCkmdGt
o+kcDeNVAido56VBkIUUDgJhOItHgmgVnSWn3zeBMcOyUhvxhQybpRjuJXwEn4La
5L/ckF/7e/0o1+jRdX7ucJB3dKXe31DAYmcSIW/1cYggsTKN80eCVGzQPHenT0hh
aai3TZ6xnxvNz17T6ULCyCCq7Yn7ogdP+BfV0si6QDp6x3Y0kT8kcSsnH3tSMQ32
RmFIVdaMZineqEslGIdFtfnU+kJZXBCqfi/QTRIxs5WJkGOeDAOv3pe3x+FEUBB3
Sz6LtuxwetYxIVpksM/ixzLVlqdTSuRMIl+BhaJir1nUMRgUUnOPk/wHj3G7QLT6
/8ZTi24zm0H81iO5DHtAh6HWZAi6F8AkRTWfpOAXTECzgtqN+bWjOpxyS+/LBUjS
R3AYUzjZ8C+D9YTLIoeTIxbcjUs1bQW9yxOaSNaU4pvBxhP00PXEPynk75gTNI+A
V4fUYZNJjg+crSumrqJVaSfavS+Y0OTcU8XaAIb+PGh74zMI3+Tn9JMirssHFkaP
MlDkEOe/OC2l5DnSQCA1ZsWKoQ5QYmYr1EkiHph3tbiKBdBBdLTDeAt64mVikRTE
HauqmmYTmWNBoNDD2cXzBcIlsODMgORMAIGbpaOZiIOONFFE+8ScjvHR0NO2DcGy
F7Q3iyyOxvvxIdeoPXaQee6bfcXpTSkoQAaN7h77wYAI3lLww4dB+mzQ3ajjl2rV
hAvctdbFxTOLQIi+S7n4y0HqN981k7HojNASEfw1eNWSb+JH/WozAw6tng/1sbZU
dL1ZrowmsgsrBiCGdUP6KHoqdH602RimU81OmRV8VRtT0J3lyjxcC+asifp/d2Be
u34Wnla5PzDmmgW3hRAIuWkZbgDrbOp+B13fegVjWC33kruLPPPC7yQoMJGdur7c
3lXQ2HlLG7Ka/ol0Iob/GU/XNohGpivJcx3J67dKsx/qAKjDxKbJQww3LBNRuz3i
tC/Ss16znVWVotP+brodJ6WaU3EAz9h2B8ltvDA1uORktw9hl5ecsXMyJeXmAg+R
LemjNUBm1RP7fCOlD0MLaoRezc+H0mN9R4EJ7rqtxdfrRuVzznw0enBZTQCFoIni
W7ALz59h5feesQU/EsiFSepNvSdOD3IjJul1dFgrUj0MQS+eC36bJz2s7G8uA1BG
iEuNMIXsBzAve5XF/kjIcK8K/NdQ9xivGuFCvmwc7wRDRO54Iit4fN9jv6BxzYAn
xh5M+MKmDkSzDSekKiJw67QY09ZFB2RiGnZqkeQ8tj/2hBkFh4wZ8Y8x5wGzVoeY
zCE/5yQWyLMhmH8Gprr1r9eQwXkf/dwQ0LR466oLT0ryCbRrqkMvIsWcLMzRLWYY
z6QaeApk/0s0ZJivwyGhVW4fABs7GAbA4/oi0bdhZQBhGrQeyLT4huSOvmoiFcoY
/PVql2nuSoUV62hMcesuRd3u0HoZwnp7pWCEiclMppanDrw0sRA4+3xP6HSrr9ZO
1s40p/141VtAWhGZHga7B/uF1KxxrZNbb9+AEX9BcaJQpNMcZfSa24TmD6+5zlAl
OBP2xPCU4rtUJala8nXUD2sH+HwktZ3SCHMWebrevEgeTGDarML7AdPdZOjui/Q7
C0EC1AfBcCR2D8LjiESfnwcB57I48KOvZADSJNlepSHM2SHFfc+4cG6u5ryfTSX7
LXc3ih4zcEgocMi00Z1l37fEP2vw5bnXz5VusVM/DFJBSgu14yYZ4a+rIRPLVZFO
mOc/Hv02vyNsVLuF53U3F7a9D7mGIYqsKQT+Hq6P899mALY3p78GdjbD3zfTSERQ
uDQRXILRMQUPkVo0iF7z4a8l/JUfaAQRxb4dtZ5krQwrdAGltBeDQCoHVwTtaWvR
b+GX6dCHdR51/AeFKudOLhCj0KkTRRKmNkMaD/7LvpkrFiGh1GqnbrM1ei11BIvD
gV0/MtIHerX5z4yqgrk7j6gejuG5RZkpU4ydoWbCh0+AXmL4uXJh0UdHtEVVMgpO
h6wcwx2qjpgRG4p2kI2ksyhqfCoG5rGd7MsFvPET9/tCM+nJnQzYORkOgUx2R2HV
FRTq9nno/WjJKiwroBIZjygzVkKSZAgHN1CM02jX/Vks2hvZc52o8qPBImff2fft
uYCX7VEzm3Vpy4sUlK+YgMuK+efFKR9ev0DyZKbcpGxnXnTW1MxI3D+7eyjcw9OE
N2OOxs0YczeN2FAI0ruqNoX23A9rRD5P+yMrtcQNKf4b/ManXaEmnlw4DHuBeccd
XjEI1jEDew3zQZgsCQs0XT22ofi2n6EqYjJEIxeyWrkVjrv4I6u9MmM6RvwypzOu
Kp/197YVsnngvZIUKj+GxcsPkpRTUIzodr7N2YswGPeQz7TEGeUk3Ja18sY0uKXK
26e/C4DJ0tcucA7y3og041yqDP5tjds4ciXPvkJOdHvCr0m7wHXpxDYxM4zhrWXT
r8wiQTbCBFs2k2rv9C2QaspMZjmjeqxfsq/C1d58tX73gUfyDy9GFVRewbjsOrdD
H5SVYO76DFIGGLlu2xqIo9yMNmCwRUq0134RZj2S/ObQd6713yEivLCLenguAdwH
5ky4/6CTG4v41jrzEBobnYhYni2LZ0nNUdsgPCPBoZ31SJYsPDs0VXfJD7Y6Zt7Y
RvgkuBfKEgrETo/2Nt4/QenRleImCXYLBk5jbSQMB5eDKDoI8rsid2vxm4ShDOu7
mARBAZxFoujMTm0nv9rU83fOa/Uwkj6GoDXJSRjYJyFu9ExA5B/SbaUuJOU72Kwm
Uoq9kmKJUahELpTmmkAEYMLPgO1GrqkDwPyq0Z/E7ZMDTGIS7hYQcOuQnfb6h4dS
aiMbWnuTLMZZdkvAcWlKQLJ2Q6riXCTSU1sdvFHP+zoKgjGABe9CwJB2+sPr1rUC
h6HacFtaQU3mH4oq0fKrbFnqIO5KyiVy6cc+0sr/2iLa4eOZI1hyjlwUs47G4rAv
0j7Gai0C6WEVGiXpQmPGUWV0rj1WjnMMHAOI2xGeW2iM61UDG+kQGBuUv1uYkQd0
u64XQUEvi0fAGwjs3GKxY40ERyQdxoyLBowXZRu3gMzmMKpdeiC6g3lOu0ig1AB0
TPY8m6RaIepGvvc7nvBqo06rQrtH57ymvzZYXKNcN6BNzXQlIuFE+I+mbl6fQSQf
MCNOeBjsdo+BNnU6aCFXW4M3DpfzMylz0GJ7s+o5BRgJ+InHJoZ1uEdEbxuRsJjU
rDBgUN5mxO89NID1og4YSOdLHQK0UPrQ/2HZu3Cm5rllKy+5XaucLMU0RfVSATUb
cOtLMZmjRulozC+869r5Q0CPanUM5Q/EBahWr8CJw2Qi3IhlwVuFXgv7cp/tvIdh
kt9TccQjMh5/HGwsP+IoOUHSz8KQH4dky2Q8CfKhuR3lpSPxRymeXimjpw6EV/AP
3luaRaKGsMj1XDIru3AeP2jivGNNhr3oj0UKF9CeSBUclyLGlyw50GDLp0lgvyp9
mVZr41m4M2qRnnSpBwK3aG5s5YgiixIf9ipcqLAkL5YMU6iPOUA4N4zQHFaLNNsQ
AUARMIUTschCZNkVveakCiex99FWC8+xgQnAl5BRxnM1zyleiuzbjDY9N3lKXAiE
/e7LIyUFSibRrc+i4/ffMV8O5ZkHXDdy0iClZYUDPnYvf3X/gjPDARI+uK8Vgd+W
QOrCsvYnN29HSuAUZsRdXknUODk3+lpbm/PYKdIQ0WYzHYcXFnBUjDfV2FLH3Ji/
VEPjWPZOXQe3SCqpkZgoAGUOGcjF/2HSiMDn56re5NoPO+dRSYHE/RJFJu0B8gt3
p4C75A9T4FI+wAPbxoXaAEPYFyHQur7O8eueQj0bHvs43J1qBgL3IfWPz3yTb8R1
OpiefHWmHeqdheIwXRr/gcN4vJvA1G8kUw7X4SQCtYR3Qp5LmY8hoi+DY4Z7VZTc
o6fGIIhyhmpKZEJBparzqGgKCmtabildyfq6qlWKw/UisZxOoOxcSoBkUzTn1yse
V0SI0ZAxBNIqBOJOxK5wnPUpmr/z8RKtCLIJguV5lSIVoIXtxSS9jubdGCFqvV79
wIxMHjCeYXsBe1S4/ChsJzWxvr8ywe3mvkWjaJJ/CibXF0qp5EKARAfH95vg2ar3
Ws/wCfpES69NI3pU8LNktKZzvh+rKMu6Uycd7zRVL+c5klq8O4VhDQooszrxpACO
JTHlzkOSZrn4mBgTT06W71NJmE7cg6yTC6sNj3SAHJ9AQlypdW++oJiaaKf2/hP2
S9TWS4m4t/JF+VQVAy7xnKmdqZEh1k4EnB4hYY6lQKA/2L0tfC9p5xqVKocfeSe7
/Ljalp16hf90apo0i5fgnoCTHhiwY96L9qRkaK5CdlTcMeMuCblhArw0giGF/2t5
x5EAtR8ukz1Gm8LGxAhPfW0/g4PAff9YvpME1g0JG12tHrcBxxiDJgv3WN0HpP9K
15IYayDh7YVTqY7GKiA55Dh911AT6A7fjSqD2IfZwB8TiURsPMFVINJSw5HubwNV
nb0yN1y7WXPkPFQWaJbiD9Xc2WT6AXM5rv0nbsqp80s3PNhk1rPpXfZtwRCYm3pu
io7U79UN52yKvvaihRxiRCgC+js6rW4JoChhwJ9fJLjudRWRVGKUcdFDH0Ay6NBO
yvh2FRiFf3AUWIkrtf4vINFb/FuzR4dKs11RC/7c24W9uKUNbhf9vjp8LfEM2Uid
haN/BHoD56zi1yWtITlC/KZ44p+q1tmHUImEaziCFqLwsSsi/y9a5MOUdmdoMXNl
EF2KIQZeZuwANCigxmWWeb8hKLqJfyn5mHCbICrqIc20cg9wjiWk434OKV1h8cMj
GxGZ05kijCKWkmewBLFy99LKHRdSXYArvObRdACvOR53/gBtkn5q8/tppJwIDeIK
FzJKaYNRr2I647TvLgHbWRYW7XMpYsnJmA2I/4SE8d96ak3Tc1+sO2atgZVZj/QT
uQL2CZMylCBpEX8yAzfyckFXyz/rSRK4/IJHReLSfeu84BG/Hp3CZiWfOO6EfMry
Zy7jYFpGG0vF1BoT8T1mfzFlwreB6ubHvrOP+snS/RIr+b+V+Z7IzGorottn/tKK
yedVvsYY1Ha8Ubm7Jk3ipod2VUFIslz8HEZxAP3egWDaAI03a6iBnxgPtH0I2cTY
HOKkkLuC76G0vrYWYfMxpFazi6+TJa0QjbUkxjCEADwQcnEgXT1iJq7DTpONguPw
G9AjaRHMStN6BBV5WIGTzTF6PL6nvth5dadXZL4WaMRPipfHHOnFMOw9s38c+qVN
PHx/RaGxtBTMbNHlzMm8blFVPmVGECQQt9jDnkObRd72XxaDSpqzzQZvShYAhmoK
56gqOf5N+4umTcvKZ/gVjut3Nluq/nTs/R9TncTIZ3Cr9xilarpXNp1+/QQAyIfM
1USk2ta1U0MUzMQYRS2P68805V1HLQwgCbkrHIBvRcJWo27ENqOqZo3MXGq1HaJp
jjUPjR5IilWz1FxzzmiVr9rout2ccmwc7yxM9tY7NmLydCsnqaSEKhhYEbqI5dIu
Tn63sBlbzBc9hURDY+ZB5ESgODakhAYz3MUNU+7HdODa+n41xTRoxzcULL5h53Y6
1jDVtnCCalg39dm/tLeFRqWV1zVluCGRdQys6e7wLjnKk2iJ3YYDjskPGYPH8XeN
SGa6WNFQ9cQpRwqgBZ1Ajp0Vid+yLWo+ghfqXMVeV1IXeOOg/IPRkqs8RjjjpsqT
g9pbZe4wc3D9fT5oIiY5I8/wyAWf5eIJVIOKs0Q+ksp/8tYiJLPN2mQqTT0B9HUI
kag8y5GEL6VCsljRrxqBYO0vJ2pAR7/tP4yCTun5J5F0QM14ACZb1NTD8QeAr/Kd
zYcSS4dFx7tGRVqqhPXv4A0YCTUEFZaib3ziFDVzW5AoWug/9lTEXvDQIsnXM8LD
24WqWjpZfhIbhC+k2fmvgyP0vLm+6z+xmz28vGVutfAFEZByNyc11zOspRbrrrM+
+jJxHbRMxEqmw77VKkvPlzxOTxNDKusS2+SOwgfAe8bM86COFFQ1FiaVKVirmQzE
Nqojad0ubdZTAORVLnuCN9JKuH2RRPgYpgX74aEDj0uQEWNWtKbaHidVpbJ+wjxr
KYGQICg1d1koVKE7K+XmkmmAdh5tznrbhMg6x2D0QkDHa3TfNcjuShbF3zbU4cAz
PdqhlDRe6gR6fd4oxbAvN3uKan2f8PUZ1Z2SzzWwQ4mggRo9O7U6WhBj3gCbpzh8
172nfNJ++616nW7pWo/dsKNzu6Gqpz6JKVtN3nD7GSF36qtZkZHJsplFclITf6Xa
5anxr4gojHrxtlaURb9/7OVEKQwsxZKIkdN651vl6PaV6vu76kEQbMepI0WP+pOM
dpN3jEVP956Fspg6o2l0Y0pKBn7l6M2bpB0U/rJ8C/wbVmcIcEILZ7l7rHPtHRIB
XShZ3Rp9YzI9h9vgmy0vYX/WU+x18inwT1v0hSyZQX21ROAuc5RZeKhhF4j3P9k0
fR0htXVouJ6E0zX9bxvvaor7ZSzZokfYOFoB9F8yQQOHLfR0XicX0o6YZxIEjUOY
tdBnbk5dxsstL4zdUQasoP53a16g3qGNS4AToHX8lwQykbzX7hAVQ316EQHjLdtt
DSdEtUhwWd/O3cIs2vl03dILfuS6JiBPrPlHiS02En9+PCcDyJ4IG2NYQcTW4q0e
jZEaMW1PDlj1jDT/HCWhzvyUw6l0mHrRZoCexp27R72mmrHvZfigGumWwm3OlvEz
D6xBsBAadvWwU14QFhh23dXLZeUSY0keBO1e66RdCZ0ISJ0+OlvxKRDMFB8OdsM2
Y6Vo8CRjqjGdjjWTf/i7OSoYhulO+z65yhfPTSzClUNSuWKVCq463R2Lf48EVKp+
5iqs9EcFDB7ouaxtxlD64pgM/sOgO75cJfhOIdqnuS2mepkbXe3WO9zoMcAKem0y
4IeAdjQWnD+VjOrb0n9jIjI3H1GAAsF+EWAygsYba2H2ok5KY44n2KXzrQA9qenN
MgG1JdAHtrf/jZLbjFkAZM9YOEqf/7mHVO4tShYiwpKHbGPy8M96scG2ooGXWmnG
bvfycIcnN/lwXVKBgtqIpWFxVdnvGjnP8WTpLOfEqQwlOa/4Ou8dzmQSIsc5Zcvi
faRZrD7zlzzAGfwJP9pBS0KfyAryZ+fn7fdnp80yM9SKtLfuMW+UFS9rrIpP5Li3
Ls7K1At3f+hCWcARei3KNH3bN8faOlgtwdxIcQku2uQU+1AhPACnX47HDQSXPWFv
Pc+knfES+lUuzsP6o0RLrTxr9qXtF0t4OZUTAT8Vz6rVZwblgfwxjS6qKGHs0nE0
PJUqDZcbFGhJnDf+EiDABhy+vS1vw4W3HhQkguuAJ9uoW1ESQH4QlTWP1y7uksAu
UQtXyFl+kvxVilJYRyP6xm7INy8quKvEhCuSWeux/UgNKSAu+VbRVJ2vqECTX0jt
3kLIOuW8gJ1+BA9L7qzBAdDQXYN4xK8YrnWFgwefft/lpoF3KSewGj+L5tXAhnpi
vj0RN7oiJJTIt83x0nZd0OBeykF0HpGw+Djf1G4C3yra61AAbimQMh3yfqAI380Y
TlGwVvipBva0GrgYweQD1a7YLV3lKWyN/brYRFvjEIpf/PmBjt9QJnVVlId2rmxP
Ak61m3QpsyboDrW7VY4V7dBxhW0e7uzUrtbMVfo65qWuWeCaEnle2EMA+16q4ksc
UrxFCCRBGlilqFDcC6/sguLUNWTH06dzdmwnzXsCXWXSCa8UKYfbHdRNDstkUQuS
vRZMU/7Iu4AbfhUO4HRjxROqFIemaTK5JcVvFmhkbAsUW+xUntxZ+5WC41IUODy+
CmlXVtbdTN8NkN+8d5F79CdQ4J7W0gaJqgQRfpIMwd5AeJ1nCohLGD3CDArHY7EK
IpRPajN0TPuYHzzHyHekRLhDCfETnZT4nYtqbOX4TugVRqFiHAUfTsKI60Sh3UVx
Z9uIy2xOPXx0b6elXERl5S+EIh+OdkNcXsbJ2NqKcZakEo1inV4Dc1UHZLBGT2F0
jrGAxMgCqgQ6CvaKyE7p41UjF8oGAUIN6m0AmJgtxWkq5S60PHqiIyBx9rRP8GeV
UyZ7svvQosE2Y7YV07M/10Za0DDfUKtfja63JlojU9aUcc9dmxIw+jGHYQB0UeK0
wPlbF8yCbK2cKmSjebUv2Y+A6sdpd/tFLZoJv/Id5QjLaj+PJboWa7QmSysvYdBh
OHdZ27SIbJed3cDO5mQ30Abecx/KZcGfWOtbBQ1vBzYaprwLOUp/zEMVI20lsPi7
ShuNv1nobazLh01qJc0HZgEA28oHeEZ6flVha2/LcDdnQnBaYAOqb01LKc4+86Yq
bClK3GF+SQG7S/nPqpcfd0Dxl9kROLLRI3/RuCBvLABSBJqtRSGTO1p94CiUjvi6
BbH44Og4wDw6bOkR0OBvYq/c4o3ZUpis/VxHWnfasgfAhCM7y6apBXMAUcqCd5RO
6R9VFTqAQXWsc6Oqg+9/JOsp2SDVqBeFv1uAWIvCkkq7/X92IWNHhFvHLTx2TJkh
1lFKEQl2GKp3vKjDjf2glOa9x2DagZD7K7WwoK9X6Llw3Q3ADvFfFd2qZCRm0Oap
EQYJI4yMVz7su+9LxkaHYakpk00Q3WPpidAXmARtIwEI3UQ7FGBqtTOEGYmqGUf2
1efp+q/rT/FpSDebaCiPzHoZ4c44g8bBAnkFP4KaOzLS/S3hVD2XIOXzRXsAqICb
ZkC46Ixt+Orrd/L4ph3CWIzNiLD5wz+tHmz/bCcZ7uEPUpGj7t42xRw/c8oK+Wxy
/JPHqqPB3XD7MlOds0ex+MWbTFMKmPdjWZX5uRaC6EMPo+NZqgYtTgdbMOKZO8Aw
/unyeQbfWJd7YB2zf21NTXBZYln2gv0KkjP+zBZ7mgOmXYyH/50cp2YTTQ71JEAg
ZvBHT3CwQj3/Z+a3r/gNEmfexLQUusPfYw21f+48dwPLHooPJVE3Z+4XXFUZrwiR
fKXqSffg8U3ka+uG0reKdOsK64vF12PUVPWvg9b+/jsmMpxskZ8zHrDxx3Q7m25q
w0XQmWb9Y97QQZt2qYh9DMhOWRM4L36SgQul0DAhkG5J5HNQygY/54KKI+j0OM9k
lPpz/TDclUo1FmktbavJ95JzqT0et7Q65AYlSlaBfe7R/qeuNyARl64E5v+OY0Zh
fxsFGtVc5D0pozfhm/y0dUKYGo8Brctf0MFdkYYI8Ot/kCdiDBVNqrAHXZmMg8Lh
b9tisPk+9sHvZEuZaSxkG0X88z8a1hvtKjMUxqXKuQamBM/nr11cvZlRMTf2s+0T
Lbd+dE5m4Okly/hF3v/k5oOlug453MgaJUvoFFMnaoglN3ZiegGVu5Bbkim4MTnm
vE/rgpnPcD65cPjDIOC71/z6ijLkfL/NIKbqSJgd1V9d8vb2O+wP75NIn66YqeaU
Av6q73y0xn0CYRChizghFdsApw5Ezu4zbtDEslswe/Z7WPB4+40zkWJ1UKkCgfIQ
Pcx2CKk7uSE9dfywgtlszBqaukvWfJ9Zs8BDo4wZLDif7QFpr3gzMK1tNx2cvqx1
qfljohJaGu1sfFWje+xuswujNZPYJOyQpvYitW6cMeG7R9W1tapTP5mV8CKToDdh
v6Ds/WqhIGkoaSDnHuRkQJVIORiahshfSY/QGnIPMu0AcB1TzhaxFgIn0GJBq3Sv
sJAal/MbGOkEGz+N5maS4suOMQHAdu1gPlB0aCfMh1SAFPXMIe4PQHbNF3+FkAFP
YaG3AUkDxSUKTo1SpcpKzvlmu/Y5RMJOZUBBasftIl3HQKr1By/hfL5r0VK3/QI4
6U45PCmcy4Z88agmtvyaSX6orQ9BLZzAVhN16Jn7Clq6QT8ky3/iBUbFo/5ad6HZ
zazoO/xnsSDplkeYuKz8OZzzAyjK8dSp8P43kKdt/rO8R8f9pAr4GyJxB1IaWOCP
Jlo32mHECV8U0cYt0Yox8Ufaoz9GpqI/9T4inQq+RQBcR+r14i4SHe5b3mUegGvD
1LhlOxC5bFQn5zkYUetHLW8t3BlzFn4BOdSgWUvFAGRWLXhFS6+NDQb2DA6lYxlI
w4hjZ40esX+7p6cQgf62giQjVEa88c9Ho6V9jYVd67n8jG05QqCdwnDly4Hvj/jI
24JD2RWTL5LlcceG3zdbu9fsVPeEU9kIzsrVVd6fWdsFpkRJiXvvDVRa12MHqNgo
59FdhJ8+/xshW4+TnToEAu78UnzHG5tnWRZD3+1ZnMXQIP20QqXzBNs1whDjdbir
b6j83NxnICsg2aQ8k8+05eXNv9ejeFhmBD+TBcrBrs9LTowRg0Mn6GSRgXupEHBJ
Ha4shQtQNoHiaMZ+Is7mq38QHklzhcDMpT3utVVmRMr2ALNwjPIwZzpgJsKW968d
Fpm4/NfSz7AuZPxp8OkutjgKQaQZblWQ87nkER5bj24Mt+6qqhd54cmH84HRXNCW
UaHGKyyfhSfvGpMMvwQ4PDV6FD5gjTSoQ/18BaPZvYbkLFKshDztwxV8SbyEFvA4
mYFLSz2R3b2QvcZj6yCUmBT/bxxpLxT9zrvdKKLpNfQX1k6jVHZyNxwt1JY4SUJq
3qTQDNDsRiCOoWpNfATO2W33hu4XRGs3y8F+57A0j7N0fNvQ3lRm7UvVF5CO4YBj
rCP9WtpDwEIqP5rf9anln7i7Bd7IRfongG8gvGnx3RuMJXEGChQ3N0RPdZiEN58W
linO4ec0/2JnxQrObV0DjIOgpZsIfRaRYL/MmxqheG9/ucsp3BwvGRiZflyaoLml
kPqHim52m1n7yN7yxTOS0kCpJ/UCAtUrReL3yDDWLsTY6k8kxkTYqive7HLxe7rF
/GhpT3/dwbw81tgBTIl1er80CyDrBfboD0uRjoIqIy1BPCYF+fwsbzyDDibhy5Ww
Uznu4DASKWZk6Rr9pMo0AA8Jq5Ygid79mWr+d8EWo28OKuHLR8E0ME/cmoANatno
NH2qDQyja5oYfBtiKE/VRFYfQGcjRMOIo9B2psTPu3HI2z3lq+S4x9vO5dSjJWiV
lvi54/vr037dEoVPuBDP23ueq/HTxwHn27VBZS03Yn1oKhDF+CpW75sgIgRf7qWc
XdiowR/kWgTEkaYFpdYuOx5IR4rqm5ik8zOAblISlLW0i8cMsdvr2iLBy5sleFDl
tcJceWY+EZijPKOEhsJjuT/yzjkx4YQLzFE7T2C7B25Ln3YHDgLhP6VfaIWwoORo
D8OFZfrO8LMTnhTLD1eV/qSqjOYcJCQx7qXXdvPCyDH06i8MoQXLL6FkPtYLIVV2
i7jFlVBH+2okmiqDkrUoJXR8pHRdhKMhnteQCgtt8ukdRlk7GKXKv8/ABTqfO7/n
SQXb/Ef4+s3MA7Hzqmi3m+WKPKjoASkUvJ2k1r3WOvicCSKc2tzWrFZ06Z+vO6Pr
4LKQRbYyTYW2mfpsPAa58KWkTe9cqvmIE7QPwCa9N+/ibH9KmxLZVwYg10sOxph6
1zEB///4pknAkAUiuuOjQCxZxaECiYF+0RBExVe9Vm/TLT7YkQIWmJaDcAQn1oYF
AfKPYrQuPk+2U8JCNLCpJbiMn0LLG53GtThU4hKMPyLf6OLIwVKjgkz6s6pQ2a2Y
Cz8qtrUtqdtlRH1Q60SSLez3dJRSOj0MyujF1qwhn0dUeljx7MvAqmcFwUCMBQ/z
XSGLtLsKONY01ifzWgFpkVXSzNnZwGLsnG5qeiTvwacg6ns17nTd1LG2jtcDC4a0
6M2cXdIl4rEK8G+nWcsi62F+DdECM8yCxFy+dpOMTU9VjCqPB8SS3k7x3QQpQOzb
T0TQUJo4AMPojRNKq5qXgs2KEtnr+pQ5C9GgUprgGo8kQLXpLZZO06ho7QyLlcuq
7CMD6LAp9ve1gXlLGhIzwV2jnCxqGkLz5olNMvl9tXDEOJPYhKdT20YCV20zYZWL
jKyryQ0gGFyGfaOx7QB7tNLk+kzNJnNnxAD8u4CI09aXt9to9eYMhp8kP8PRc3/s
sF0j+FUGqFlwE6GvTNHm/lscY8qhTbBmQFpXnCN0/tAghu2Ayhk0TVNrTpizM1Hf
fEOoiw/dbIepkFGtm/lo+uW5VrJYdwNO6SHU0I+SL2GlTZeUpenLotQlkQWinW4v
UWeu1SbwEGIxNrjMi4xhzGYv/XlF8/V6rFbor5UbPf3iOHtMJ+Tmyi67agDjUCz7
RXQrbDSJnpcai4dF5BDsKy93glmtgzsauRORNv4xoRKOVbxDoJpUiRhzj5X+OZ7H
4zu+q4l3qENCH/fNBIe2EGj4V48kMDF5HkIbhVLwXOXhokO25DUjcNemVIN8eBoR
teW0RfXdOfsOHTWLZ/5NqqYcuxloSsdYCRZMhE1jp2nsZINcvrZe9NxG29DB6dFD
GkJKudlrZ9yLgi2dHHm80+1p3iy8NIsAl36hwOJl+GgaXjPX6sShRHyst9gdzJLU
QWVCn5+UjS1pITBnJ43nVk38YAeorAZozxrjC3zeqP0pU2Kj+HkrgVbS+PywmIfp
CrxJIiZP7jfuoXG/v2nN8Au1qYsWImAdUuzkosyXLn5ZZYi01BlnogA4e2x+cIIh
ZmvVev+obRmf00OUjP1iQ0JXntNfMlBh6dWpcfmTEpVu3QlcwF6dunf1S/RG3vEd
fqLl5n6+ZSNTt4u0sEEl/mxvgmOuRzUGtNNACxtqMEF+XHGbrTxn1KW551kfFpC2
IAmJmvWq/+zTtZUYnPb5CiJ+HTr3pvs/gVM48wCNww/deBj6XT8LEwz92iku7uYQ
wxIaLDEuf8hRf3/1wxQNLFpFnpYa5g6JePmdpbfYy9aBQb02yttADl+UlNi7II/1
jR1dzzgL2jHPPV1UXfbOpbS2hrHu8tgA2BEvnYtDHhhKjo3fD/r3lHKaTNOwISNg
rzugPd7ylz+Rw0RZH00g3+SrIfsTqsZZ1De6PAs9YD4X8qdlOqRRKQGHisvu7eRU
Pi2/Eh1pOgOXBzqGK2l7JgzKT6sxwZZI/+FKefjvjzLFB9sdw65UaaC1ElgpXk3J
/ZPbthRzze84EXGKxcLw2s2h/N83s8dqzt3NOwRhd2aZQvlItXvr/UerjWWH8jtR
Gi3R1SdMj2/uZSOlz6L1+9rY2yMYzXuyQ+6Y5Pr7LT5f8Vn2FNKfPFfO8yYJVKLy
tOA5Azy0GniQ9HV6VgG4Hi15Mudmz5hk8hvPZ1zdTQf7xrnCuGRSW18HcaTgJUMV
7ZzvAkPMZq8RZ6iuso5Hd42GiqbQO4sC9/5XdM7aqlPDEZFXDMw8JQGKPCUgtBEK
YtgQyCUao/rRix79tLHSMV7qOZdABLerb57vsB2O7jlTC4YInK+nTK9tfcoNFxnG
5mdf2xDtn1izqF6dGIlmBZsN2cqaRAIR6yaBv0s/jmgpFxmE8ted6gZ0Y0iQxgOS
/DOxE5P5pu6rkm0ptlDaCIcr8CjDuJ5oMWAstEeFaiiLUQQaezhml99+9MCCj2DM
0pvwNglSS4GWOVGI1fXh5t/+fKnMz2aWcnVUKi6l1Jue2esvAGZbSCzrTNKTwfHU
Sna8mp0oZMPlUmYCMGOgguIr+QZq3xEfnKdC4FGbvftG9YGuaYikR0n3xZqm1f+S
TSe8/sbMdHc7vMb4ZfEJwQV8gittcjMesi1jGXgfwsOWH9X8VgZHmTHFS+CPfOmU
knnbjjE4Yt1a0MJDszC526fMm/a9Yw0gYjsTluf7kuHgg84MNGHzFUUuZED8w9Z2
bO82FK/Yk5+kZWBW6txa0kEF1vlmOuJhm0dplSFMwGinEQnPuCP9RA4JJLKNsAH7
N235oaj1j+7hV7eFAvd6OzIhyAtUvoDFj0W2o8oBHfLFS9UGRoJ04OPiwjbXCMON
LNiohA5VY0IyWF+lwL2UKiOO3wK/PRJXVLy9TolbWV2iJnZk+OqgHJz/qu2u6RU8
FMNp9LskXv6sRBPw3K6gSwPEVAAP5am7peHPTA6Uzscxl86KIwDaoSignJ96jsNJ
E9sPcRR21xC8i6mmq77EuwpvrJwhyn47huGmcKaZImoOLYWr5dTbN5kJOLOJnxAn
txIckXqi7J0r4imb25rurG0+FfuIe6oCnCDI9Z99qPaMCApBoCH5zVLrTITmjdOz
Pk2tqmmF4jiq7XTuGEzbziSckR7jCbTsCME9O+gNGJGiHNzanbY075I0EaWztE5E
3eG+P1iinXKOuroRUehkoeOLvlY70kuGrgaSQY20Ch/KidTZVdghmXBZPxRQqi1z
rgjtOKMlzp9FhJMmQGzX46gGZ8V6pH+A4JfjGMsPsgnkNINEpdOcKmCE7KI0fZAb
L1WNsvqmw03V/qUAjRkn7CEy5TYfJKboj7/IDtDojEOFnwtO7x9VdgDXkcIiaFfO
RWrhxb23E2yQCrys4EKMTe2cIzeMWQy5Cw8YzbyzaZAgVhhRzgXyj93EogFcDDOA
y52cfym7LcDNukOfiDxXn/G70MBiP5vvmJzBB5tEIRPx1Hz8ul/jZqVs/jIJFV6L
D5Q5JfvEXob9Vy1k0ePlNQ5TuEZA7vOqEpqe1nm7jdtX4jT3ZVELWLQg97qNyybd
VT2vshn9VEBsnYSlkuJGYm0C/nI3i59Qjm08C7RwccSqQzU77fY+CVfel46X5qbN
qaocTYcjupdiIOWMuYbmilB/JD5eM6s/TLC3qiHekEg98JjoRk/WVvwXxFYHJWq3
39JyhmpaHteNNHwoPFMkZZC4tbrxnZ3/Mjp23sOcfOjOfyE9dXtUAAytItb0Hr2m
5+sF+5fUrCG//hZycF3Tt+RRy8kfQtV2khyNLPoRo5fxnsiKlEa1/9Li+FvJrzem
FyRAwIjzSTVxdElbMz7rsM5WMaVHb1BjedGGYiPXExFDVTVH0AkUB3auxZjsAw8t
TaRlALudEz6PxuTBjhHZkbluhXI2+0TpnHBQ/AK/PA7U6D50yCN9LcRvubjwdMOp
DdnnmeD6zUsh05nHY6/ohPQmE5EvaIpZ+JxFNatI63P3ltvkmSfDeBeMIqVUPZbM
bHSxzD3VV+P9EqMkeeNHq3r6HlLKkqJPasx6nsNAizlYcztbxUzcYh7b9bD5o3cm
BOEEcob+620AGaFp38YsX6fJD7dW8mOIRZ56AIg9D5BgMw/aQ6bYMBIWpWO/yB65
XvYyH3+xpAwHU3mLjjee4moqAqTi+7xTBeIaIMh84mowEbS+PfpYqOLKAEPPOLfA
UOPXYjEcd6ULSGo6Tib2StDQmwY3uefUjlTLXNqVEVG/xrGzlImJaEmNnldrZZdI
dPuQ8Opj8LsQQnr422PCVk+0JUfzd3KUsA9FdLzoqWa5I/Juc5dE6GdBXUsP7JSf
6gRrw2816XjV9jOkxfKnTM52VY+bYD+I7yL5iu3I5P5857Dms0/4Q5qOEEyZjaRr
UopcN7jXHlK3du1ddjtVSvFhjKS5bsya/N3l0N5VwD25/w7xwd0EPNNp3k2uNg7v
IpUcCsY0M+pUqTVtHayNLN491KBBKGXzUW40h4bSrikqtp++quh6Klga5zoXT7mL
Q0Jcb9lJ3gO7kzo4/0C17M5vQe38IhKN7XKR2pQqfQVNGrCT4WvRB0vhuej6GQJs
ag2oTYPOH5p7eq/7h6obvYPBGEpdc2Yk1+/hFEf9goU+bk5wNIHFfEfljY0/ag6d
uXk/y77wbbQKFWMuH25aUxKASwNXw1dgwtod6jt/4AXCUmai4YXpNhtCA07xH+Yp
fE7zGcku0Oil5fPE8+PzJYbcd82+EWUp2lowlYLL0Gf5zIfYGskASMxqMncf5Wyc
DOBI/QKhwPTFK+UY6j6I83jFx/T+DBUuqtWXfA/OaK1Uzsb1nrdXf+fHwYOGyUDS
4PkkusrVXseStyOCALxxu8Qo9OA0o1xm9FmuDz2n1jRRX/OZBpxRjJQ3wJw4btdp
noyTBmuL6Jfhi9NXq2R/r+InZ0j9bznszPMmw5psNaTY3h87N4K13zpNgEAoqCqA
jknxmtEqB9j2tdUrkIS7kHpBPfnO0uxGwmEWOYa0WVBDqMAdg2V8ttvIFUxgPrS9
XTLnLBY7G8FOPgM+XWtIDQAV8Nihj/kut+cK2vQaG7RabVjrKUIjxUqk3Re77VGu
nLdw00g5zPvQA5uAma2Jthm066HTnVEjt8YIzmS3O13YlaqMnJEHyX2cMq/gqWNg
8My6YU93hcd6r9au4U+l3iYcfEvS9rt3kXPx+IzIgVXTkBCBGb0ZMgfyaxRZQ+r9
eebohXEm4jnBDL8IPIuAH+q7wUgv7nySK3WfE9XvPQ7LzAIiUXvsEn1OLn6l03+I
8HU3vTXcppipFukjG76sHCnDMYSNl/Eui/KtSnh0dcPMg7kiwE0SBFsq0hMeEEO6
savEBOdtobpEBmLZfmQoiLJLOdYEjE6CDJJVgCUUVDiUH7TSHaUoxJ6d2JK2oACI
vrxKbple+QZbPMTKyYsILTu2Wo6GXfNphucX63AhnenprqTLFaAMSzOZk3Fgv4c0
DzKXbE5nDCDW4KqfBnBTiiq5tEiLPS+zkvcKU7YIaOVi9O+EL7zc5Go2iQkU1nHH
o0aDB7SRhGXzl+tzDgbtoEMdRCpvTx7DG+y98s8b/KYDl3K8IfaqZkG3RsqIkOsz
men8yIyYNLlx1PuzC8ZcbtsGJTnYJYaR49tRI+AZnCCo9bydY5ONveh3H2X/HQwr
JCjyxo/W0/kHum58HkHoRZowl9p98e/NDC+Tt+bgpTtAQ4EBv/c/BZSpRM3XuyJg
xb7tHKXJNOG+bA6WyG3KL5q978RmSNsYKRFYACGie6OpOADzfST5e7Ykz4BjqV28
9KIUKbVf5m5+JhNcyvRFf/UrgmnEvn/hz43xb6yC7oXhLKqcwfcgM3lE58BI0SJJ
14Ab3Qg8cVR5z7gNBia5DyZnkyrK01798unJGnfD2GoW2T9V+PRJyX/jpaDjG5Vj
n2eE5k+1z6nl8Z3KZBXxep/mIfFQOtPQHrCMdPO9/+gTGrPr2Nthjxuf85PUFiTA
6jyhQ4ZhCjGbD4qzsj+BMg9YJFcj6pyDSscots02cgvo0Fen31yQODEHHeOlaG2s
4DxRE3FXpzKdvl+nYOtPEACvHkzv98MWUR0pE7egX5OOLC9ZB1OYDWQ1U8ZVTlEG
8pxt38M4d9Dqv30Ak0B73eCaDUZh8nsAhKj6HF3AQcmkf6giAWQzUXW3JbSJDtvj
XnS3qHJxEWffx6Lr8x+DZsb7BftpaAKBN8t5AkUY/ekctqzyp0L46aT1CpGFzDG7
pQE7+dN4rQUg5336elsLzirLGV6dPRB6NHiNhrdsr7yGINyM83GwnduCcZYLcbcg
D34xvPWiWkr7j2XUFLmFDMprEJTBWElQHRAmAJMZXr+dLHuPuyYcwj/LOHMevE8N
SkAPRbeNJRtFq9ZAkcJe+hnRWOpF2VX9msrd9opfdMy6lSjgXLl2EKDXZX92hUzd
jkWrZUlj/Vq0oH8zDLkhPrqq7skA8sBPVU20nCZjRoduVpO/l1VrJdipCoxLc6n2
1FibPxUWmurjLYkOV4lsILtvmWYwxViisWIB2Ll9LUZonIwDY3NGO9h6/aX6bOA/
NXNKb8PXHYXl/ZN6rq5NmkccWkOCXyjrSZa41W/lzd0z0P6jT+0oWSeE5De7RZzJ
a1ZTeihmGiPKzYMFTXim7+a13Tpf3JLn0SkkdQYPpJ9t0gag59DijasV668f0o54
8DLSC3nW0hx/HIWB0AZSW0ad53NOQDyudq1t2OB2mfy6p+kj/phQGfEw3Iet+6oZ
D1to0HBQW/z30etVQu+v3F3gZmVCBcRuoElV/FDlh8ELyohFoqmiqiQz7csOsc3u
aBldUM5xZ2d4FhNpHkUKayZeIBTE5o0v3Asy3o2VqnTI0Kyvub43pe4jTdqMouuz
wgufWoW1OFG3n95I8HHtZQgj8tH/C/Q8kPIBH/HI8bwSjJldz1mKQrhT/RPe0k3D
ylipIlhSVFluLg0HQivHu/su4N0Gi53vQOYc8Un8ilMsol8yEgb+3Xhz1BxuvGFX
4sXm63LbMpLlzhuFKsvtERjvDh4dJ99kiDieyJq3pQGzBn4L1IkjrxoZ7qoH4WVR
ZiO+rVZxIM6o6h3yQcidZRj9h+2J1j4oJ35bJ+KdKldkNZWUzVbS+B9HPRIghh5c
zTN9yjcrudq14s959/+7tSo71894jdjBkgIRE5Cfs5w38YVs1VYBo6zmnp/eodz0
CjVz/3qtWc1xZwPi372totN8gOJvzScjiLko5ERSIKpeR9/5KWKGnTo6Vc7HNVmp
XxQsEBMkER3vTHb//8s50GKptua0Ix/g7oAxCBmzmfS8LTRONkPYPw66uFH1UgMV
Fy3auQbclHnwFt/osAe/QnpEzDI8xGZZBJzeSO3RQGF3Q9nCsFUXkCZHnWq7qBR/
EwdnadhprUvx1awubq4KseFu+l2ujaJJMKoclc2ox+qjwU7Em60mR6+IMP6aO4wo
r6S2POD2UjWbbD1GeA2TMLwt3/FWG+IuQCP7nJDJY5W2RMy1TlEM9N9Co1L/16qr
38SF/AKeowJ3k+QyEdR0PpO/EYE+KJHmwsokfhmzceS9CCfPKVQ2bySCbRA791Hb
rJLaTQTaq5O2Z4Jgp11g23WtvKa7Mnxn2DiVWWBvSmWPkd2fpYko3bOrKrxlTa+Q
NdZPltVryEOTfoh0Ud9IYfei5PyJ3w7hnfwhimnBbODKh/faIZJOTrrQ4EJIKI9a
uUC2ER6sCKLWK3rB9usej6rsUyxNFKI4LFZiFE6gFF3Df/BtwVQWh4ERiG53IXae
0o39ZoBpdN/6uYt9WDW9AEEaL8EQICA/z1Kjba4sp5UhT7KEhXzy+L+sYQoHMo4p
zhj4waOObZfly7zhP/XjwZQ9xYOdEq8/G+tog8lsgsD3d8a2Jc3MZ9uhcG7giery
A81KEgnmYbvpTeD5e4LJKdRZVn3zMmJkBkrOQxsXyfFibIgwfBoOLFw05tiu8nn3
0mTOAdZiVLtkw3b6fRRp5qI9V1UBNq52d9Anh3cnwFQ3re3RnIVGbMCmjz+BtWfN
ciPzxPzQdXTuSTGVc84wRzhsxabWqmjHdpxRbfb9SpsrI0Ne4U5ImFK8oyx4uE3r
sF6KNtFWvHx5IdMqMEuuL9FnQvw/VyCwcr6ChAy4Ug/BVWQZZ3O1CQVZigBt5QdV
y/eo15R+G3LHTO1t2Uev95KuKxh7DHfdOGoxbxprUv7E1xzPIyCxnqtZWwJUfPPB
gGSSrZW0xgzQvQoIG2Enkn+H/aowm7yWPO6Zldiyqhe2+PPZL6aEG+IK3olAQeYA
aVDPbOd68M1TIetbr0VRM4Wrn6DcnGv7AsAxPNQdOFabS98jntdhw4y2Neb5JZbe
8EEdjVylTwcAzPLW7AZ4gat3iwZusi1lZtnOmBipFVOlSKWK79MWOjhhTfYEru/S
tq6pjQFAVpsBoLDFKr11XjP3kulYqBp5diyym4RRKhgUldTxOb5WP1FWmbyh1tXt
Hgo/+SRv+ekD2jYv7QMkAmPnDwDE7T5Hina/Jv/dnDyQNIx8fba09FCkZ+/BWjo/
lC34vHfEpXrPz3sMaAygsGLb7V1nCU2SO/EBdKyv4RX3z3d5wi4u+FPUSZ/INtS0
kxJ+w7/M/y4LGCnzTLhV5aA5PBQemrIp+lx3InV1x2Z6slIL0C8FBhV6iy63vMkH
7lNSZ9cRMxqXfGw9qwcvRrkXMTQ9LArgFiadpFeB//HMgmyv1k4lHbVDThUEk2kV
WNe6SAJ3Mnac+DIfps0FTU/HFcGf7O2Lhl6VwVxaYawvow51EWpVw9mheey88Vm4
QC28xnCCa9q6OX7bhaoyr6c+UQF1xHYcyyCs/jBXpsYSibgSxQ33YOHNbeVmEHtf
8O/xncl534P20Y9MMIWLpWrzGGTgAYlqUsEtTMPnsy47M9ABgr8GtWe+NGCFumRW
BWtCIZv34w119mUgq4UzUP26zNdQUx67p2MyZMzaWdt7B2CzjwuG9nZxi7NnHLe3
0pjCO0dJKs4fYC4/2y6I37o602ipEcSBp+NZKJB5xpQG6Pr86sBrl75qtF56i07c
7icmSSV8KtBnbkt3pUMA1AfoHvJSIsjQAQaNN6+Bu4YHYTxxI+hpTDrvzpwEbqXr
mx6gIvhQ9mWS/KAHxwYFcTcXIv8rfUOn6ZzJk4AiwoAIU/6GE21bu/ur3BYLpwnT
sVsDJ+jESve6bKGqJKnNM3jDAICXMpQNU9n/XHVFTlQzq2Z9Lj4hVZ84AShmaWk6
JkBRuYUB1yZnZq/uhmfluezIYmbTMc3jNFg6SXJLJCOYC3fwvdnVibsv5vlhcWgb
07JEOciX+qIZP5YFxfJ+Se0xkNytGatshQYW0XDrYAGCbxFcJTZtupPrZ5R/7C/Q
lzpdARNaJeA3ygueW9aN03Jgdp4VFBC68XWry7T50qZqsWbi9SFi0BpqE28ojDa5
QzDqaZdoQSF1NWzePBUf00yZjH6sGo5qW5KIGHWSqFjdE1BeaixlhzTPkhaOZPp7
/DPCShvJV+za7tKZiqJbWhHaz5E/Uep+v+bY+aOCxKLqhp9xxObEnDvzi6GV9QNk
Nfw0YVOX/W16F0eRJ2V0AVLWCsJnY4EQo5yG5gUhU+2qps/HLgVKfMlFu+lh0Exy
pDpFIEMqPgwbhtY3h+njiHlBX/MoGqEX4szjHWR46R2MzPYBgeKCkjnq8QSRxZQ2
TAoq+gAmgjsfgo4BZNNuxG95lMWgSwAuC6ZvyVHul9NsJ+SlY10/ual3+xIiw8ok
NYwA4Pg9zhPppwMetVBoaRe6tgpQ4KWDFFx+f4ej5VUW0waAINSikR43MJtqHAVX
2wDjGTuZMadN6dXe33u11CkwBKuO13U2NcsUcsD4XiE5k3bm/wc87kjZ0/qWjaF9
IjDyYv7xfv03zNS1K3YZ+/DyWN3IHNibu0mPyVwmnl/g9pTO8l571gsRqCjuUGIJ
xyKBzA4ngst9iVcCeKsaQZfHyssCysYkWqMsUYob0F7Qwd4ADcHxffnIVT2ZqJ2v
43uLoWfwT2EDW+UXx1XcD/iFjkDhqKPflfWiSm0kOSyk5hqjo1d5uDNIW8psRtrg
m1tiir2oJArWMQlrF0hYQA/dEQQ0XKmMK8Fk08xK4cvJkJ1cbOqqV0t0aOx6SmzL
+DWwhWnDnf1IdCybCCR0KTqws6hSZJpAROMJWI8E6KnZsMIPXgzEgxiYUfvKntXH
fvjt54iZXsbSG9t4XPpNZLHmlqlDCgToMtmQJMq2VA/tDrv7iDzJ3oHnCcRJAba0
uS0Rokqq331wk5yRBHuss55QsuldeaXrQayXAmmHjfnw7dyc3YpnGElgMPPcB4Pq
lj8Hd/+eBh7+YHq90KbPVuUwKytOpuERaz4dab5hP5Hrks6g/EDss+nZhPDl8xZo
GBFTWN5fPr5tnQ9PZ69naCrdPOAwpH0/l5oCJlJHBvxG8JpOqkyS40V5MVqnHF7m
7luJUyoCwc3fnyDujYoetatM1TxmQIBY4/FLUuAm+Ea/vfSXlcJhjlSMgqhPl/vs
0KjS51Ybl4WbcfIYD8UubwaeDQ47HC2OG3Th6u4MfN0iBvLpa9Hgzulhi0l3NUUF
kiqOqRuGiDNZiY6f5k5IbWEawns7SfJiz36sPubHd0IIbrGFGOB72riqrOZSJ1OA
XLEzlkVs4odgX8MFqy+wEBQQkbvtTOCyb1moRix8yHU98ma/hBLyxoBn2xIOedjP
kirg7pvNgJ9Bm8CRv9rR71O7epuW2uhJhVMIl3aP1PGUrChiIj0vt4bMp95VJCxe
byV2NFe2rZTccVvRtKJWyPsb66tvRbW90zy7GDQwlYCwLa40L3HoL4hRjj8dJnOb
kkcra2Fc0Gz2q2qgJBRJUuWhmSRuZO5W721VmaRUcQwAQEwvz6T1rDNzXrkPr0r/
fV+pm62g83SgyDsUp3bpWXUYT97qLnsjqxOLmmi+BzxZa7vB1Y23HZgHRQyNwh0X
IPEJQLpKN6fxUiu0qP3Pmb6rTktGIptjeuLnAhEwpf0CLphOqMKK7PBXHDekTzuv
o3lksOAAIALlk+kcWjI4AlCXc0KKAfawLDK7doMHPrwFfPQAj8qC57Ie3Z+mdm9o
6Klqp0cMGYC8N36t1RX3Jy+WxSLebewVntS3Fa7enDwbDaeOXnKGDFyBpZN96yK7
fjZNd04Exggp0eiy5bjkaL7gRvQwB2HtCZFTyyMycs1Wr9FoPP9Mk6ZWKvdlxkP5
iaTb+eCU38FVZN8BhCiNuY6/54Ochpx+eo/MFg/6TFr64Q9rRwo2YlP+p5SWAXie
bSlKWF/4JWK7JLnSM80ukAO91hyUZgRKWokJPHB/OTppa1M8Nw7d0BnQLWZQC7Tw
+EWJzxXXjYRn0s+mIOldh0nFvhxqoBqVbYKii5hvm2+aqEHTC2rXteuba5JO7wm0
tj4S9V3M0AYSLt13MooH4Ypz85tjoCbC4GqGEbReJZ4zgodtDLAc/SHarfl/B2jC
QHHTX7OcaBMbY35EHDiO1G468FVy/ZR4zDYfBKTuSYszszkEmZ/Fjn68W0cFTTu3
3l/tNxWpwGv+nZQwoI5WK3lV3PIrPu2KvFXPiHpSuWEDI71/STJbJbuW4gP1Y8Pq
HWxGGBjjk+dafsrIQk+gNhJ/AfvlcZZHb7t8Pyw7+wePI1WX/h/o7xO5k2+jyJes
z+Pbvqoe1ahGdXHXJMYda1Pguz8QCKt9lAy7bYBNyK8UbrSrLmF6AHxpmjskRawF
S11rDaAuMcJHqNNi+R2ZTIqIxoIF+CTAhRWGZ+0VibewarzgtWQe4/N0KqrtMlaA
B3FSq0BIbuVCRoAapNVSsqBmll0YC2xInhem1JZlcwmzcY/nlJ2Y7VrWmjyK1yec
miGoxI/Set83q0RoFm6LCDb73KQ2KENnfgNN456r9wynRJDjvjwDn35oHvfpjSYv
jBJVJgzuXwaTcEpDge77tmeo3zjThM9/zbAtYuS8oCO7SrqYJC/o7WJ2TJHQ33+1
+u85s9oAJJeDe9TdLKRRYoqKaI11EXh0c7hfvxSqjdG16zC2O7gO1pp4SrDqpz8B
5yeddEsxG+XmTjv0ndvlNJbVVH2lg5ERa+5j40oodsVDDVS5Ve9j+8XQ6/uXo882
YPZaEHSH49WUT248f8RpSFPJCid0RgEi1po/6VGlXnYb9J5i3gKMCkxsfMQkKBQB
CoE52lNY+Acq89n38wc1rm2agOhHVVzM8PD5ELSp6xywlHTFbsnFVKyXTOKHrgtC
JO9R239uKcp+ugqCRGaBmR/JVKlHmct6ZUX4xYL/HPwgYDOEGRb7ZOLEOiUErwxM
mbKQg7/CGiRBROvrAwzID2f6RIC83+O9jrvQHU+pm4SZRI8xKe4ioEgxbxTwFaQl
sPzc7PsEpc4JmJLORlcMbHm+XszvMYlgYpvmr55aiYBCEOlDvgPFuAyU716feVrs
ineXHR7SNBppqJUc/h0ll9WWUQnV/0Zxgp8rgLnyqRzDI3e5oiZ7gazAqes4YLmc
2W6evnjIqLvyghCiu59SuRgqAwAekM716FaeVu33ESF0IF/AiqCWPTGF8WbC2yPW
w7ZsYxCVciT3iBwTig3D884FoOPumPjdfssaIOSirsllILSMTr1ZubowUL/bbfFh
IwtZ68X51IePTr4ay7GZR3jGc919ww4fLULSoFrOvRn2BE+njVyFYgMV7hFW0DS9
4m1bMqybSARMFTiUmbLxyy3+awnckSvUToXMQVGMNnlx7ZzUiw9h+R/2V4niPkk1
4ZrnrdN2/N7xgU041BFEykKErFxECqSEir0ZQSa427cxLFBLteBM2QFB96QvhG0J
u7/fEGOTUDe1E+xn2HK+C0DsLZwL+Lgm6yMcv9zu+gn9JS9efwtHoxq3lfq7vB9M
3ZMnhU5aI1EAjPNGyKAuPxrVUbWWMx2ODSKZ5AqJ1EgFxeWTLFViUvQnNcLTo+Ji
wKCuEF0wWWys/t9i2ThWx/+zGVIbJP3urTWqFQRwKKDGHQNyqYkPnjYvuwLf+tSu
6qZXsnqwySjhnajJ0ZrgpJ0C0bFqN4ogyQ8QUKkaZZ0GuuXwFT5qOUyrRBgxP5Bm
Jswakzm/4UC/EXrRqUv1c9FZrS5cEF1/IGkw4CorGwBZ9jWvT7yvUWXLubea0UgQ
5JdmS06flSxAI+7qUup9Ps487xZx2jtk1iQBYn3DznLv1qcKOKiS+Pj/l7Kck6rT
Vhk+etwHQOnShzXH8NIe25jMjp0B4MOYlgplZHD5bOwCE/5IYkJn3NhVnDw5DTrA
pDDCn66HN2s7wX9LaAghbW9IGVJtP2RifWm46j0/9nQ5LnHGXuLp5WsTKgxg7KNl
0XUD/SGTsal0gR8uVAS7Rbq+GlsULmxGEs7ntygzgG4SDuSGUrBoE0VBBVqkqKX5
HXmNjtGla1vEBRFBAHn6oU6RfltDNuAfhzNjWfnTXsu8MmOT61VPqwrVJTA0fQjo
rfRIHfMeiQ4tJhM9+peaN9h0KqCK5Uv/dr8ED9LXiwki81fS5B/dKwmlTWxnqmSR
M6a1kDLRU6OAdiXKXa6vl2/yer8citOHUJ43zCAFOdoeuQosI2mmlr68zaKtbUGI
vMtdBQVa53qEZvs+f4LCSQbc7CU/hXJPSJ8Gm05tRpvkok67KUBnMxWGoHAwquZq
W9YgAhOeZ9c/eXGjXzWMcXG6H+P6AABFURmbp8eyu5bR3GjWq/8wWLU4jqAESoxj
0WcIKZGwRt0p9JJHGLmM6WRWRk76V0vefQb9NmcQVVykkhLuyfiF1kDlyKMjKZLl
0abRsM1mnhhCHcVTwnsDoEPUeu0mTntYhSEuSUt/ExW8DnwzguB22N11/6kHfcV/
rGhFCbm1hGOFnJycPRLsvsWKUz3RDldiSBwjQAFv8gnOORBOqICskRoNAJM6vxpy
c94XTr6qZ0SKhHW0hQhF7MAqQpxvJ6FCxVQ/VOeJFhfx3rJ4jOPIV8FjnYHerk2N
8r0B3WPTHIoAexiP9dcS/W6wJXbx4VAS6M4snELRdu13vyAarqrt/rxCFTC5UXB/
5LxqfSXqcE/5TBOxzDI4FyNDzOB+Fduf3u2QVTIbWDnW3JebaFOvZT+2Rr7/QxHn
jVGVCWVMJ7WPBjRM0Y5vb5IkhrDpD0PRy5VCO9JGzqqKpMztb3ptYWtMTwyALV2V
1U6FQhfHamR4BfMdSIHNln3JWF1CLSfsdQBP/m/PHf9R9GKHvbwVnin4PBwmzrLg
t5bGHmUAvr9e/CvsNzPPcXBae5kxbLB24rA21o/qQmrt+Kt9z8+TqqhXTKI2Lc+s
5slo6hU5O++vJ+tGonfOwZ2cX7naeDguRFF83mAZjgBB3DkP2FPIUGj2NPXhvmEU
x66nv+mYIURpxONPofJUBi+tgzYSCNN1n2LIOHzA56RU6nRE7JkNMWDX/GEPIPDN
eBPiK8SIrH2KxxWykemXmnz0EiYV1TCpMC06SOaW/Ld3awZBU+WnzFgt9OGdaote
KWy8v7vTwDH2lWu50xFnLIDi1QUyLJ/xCo4TQe2HVQCFdmlHvCI2VozJNYfkPwbI
i2ApVTunvym07jftPK2Zt+3bEYcJEE95abmy6yv6dvoE/aVIuEiJsHlzoKFj835W
75gEXAqtav5sCvvFTW2C1poaJYrpEePdV9cFZi/S0lh4adl/EAYlgY7p7+haDtXS
wlPm9GMt9hYh+sGKFkj3accIxmcVgqb/9egQpwAnyGO5Kmz1Fl6SYLSdcdyOiYVi
V6TklfmuJyiy/aqUP3UgQBMf9ANVXPXHCQ4pignDBf1+6t7ZvCWSZaX3Z/P5fbME
54yTtRmNpT2rvnWqQS4Jp1ZCGuMxKxE+46fyvdQfdjRKj8btdwiuYEeT6eNK2gzJ
r52O3Y58D4AocVQ51DzUxKmLxvxoYCcgk3oV5YZlLpSe4q1qavGrVi8PB7yGwImV
3BXLkkbBSYVicT8HgTJzeJGL9XLtkofaDZPXGLwvjbp67GF7gT4DZn+MNVAWSK+q
d6ibwaOxHKuxybBtaz/suDddc0ZqrA4VviyHskJ/hbCI4Dpl/FDIR9GVGwr5+lOr
IwLtl0q+MTwn3SJUpC1BXbq9Yal4CA9J/KBCyPwNVQrwYNqg8w/AgBvpRVNWSKwj
/38Ds1gwJkxQx65JMQFqM661b3CyF/iO+3VwTOujCqrDtjBD6a3URgyGZaVDpC4/
7l8/Aid7HQOen4XaEULbPVs/Wx+aaBO5TeUXU0zg3EDclvw5APxyZl45NEi9W8qZ
NlaSEP1BP2FKrbSogUNh1W/Hu4WVJyv94xfkOvf7IJPE8sflGoYnkjIDeJjFKEJi
BZYGVfeA8+SVpDH4WfZaWjA05bYJNQwmVkXAKU4KbXJMrn/JnaU2JEIwTDGVY8Jh
WEPB5zp/BlSnAuOXVg4MihCjtAhly237xFQHRXZXzM0zpqiwbFk6/wCPyf5OKgDk
nhZsu1QgIpOLGJWgrGRGFWHxAqUF/KLj8WBNltjBBn8ZtxeAeNv0gc3hw0eZPIO6
yo0q85znEpCLn6FjY8TBq2OJvr79iRSCrMRc/fM+AgDgtOQihT4EnlYdVP5jeEGK
APkugJ8vDhwg73ZHfgbF55Hrs3o2PhdypEJCLKBbcbweQgp+SXYePOwVkqbPAEtU
2PKuKlYN5wE41krnEeVNIdRxMOU2KnMrMm4q0Rir8/ggbqTBT+Mr14C7GOjNhvx2
Ci38kg6LqfAiYkxIjh4pepoQCJZ65Dzx/juDqjQuXUzMra3ic4xTrbUV9mTfVc0G
MYw5FJ3+AsLYlp4icCJ0J69dnN7Xmer54QU0H3wsZxscJar1MdQPr3g5TIyon9kp
7oemmkpraAd9azXVKBfTw/BQuoup+inewaO67OY1pO6JXG8Nt0OMEwH2uHchG+N8
hKX+8tF4lP8iVOmzt9nggye/Ten8yR8Yqucj72CC9TR/SWpH68Mn7y/QwhE+J0BX
b5iAwNPPy2ZW02nqVhbQXgehzBKohR98PUnhJ6TsOUIQBPhHqrKiCPargXXOLftV
83FRdCHo+gC5xOed26oPqTbSGWR+fUhPBYAU1kBjCnjoK3UFQECSdyxZOEU+Ygbd
vbcbLv0ibNJTHhgUQbxGfcxXQerKdq9iP36j3nqY4BLDHIkymQIvmjhN8o+lXRKi
jFvamrHBuPeC1V7AYDVMyz1/7BTjMHLOKnD41KiJvRM4bt3gmDDSU7WqbTYvuKwA
GBN/n1RVrVgsR9Z8+3QYYvnGKGYkybKaseDcaffX2yn/RHGO0N6Dn69dNbKGLnMe
cdjiWLqgoHLtwSo1PyFqqwCTMYOy+lakjEEWwa47N2AE8iI215bPQr04qT7ILKu0
Sd88JHF/deBetAWbwkrqwTOFeXIag/Neac8OH9fAJmEglG+1wV+c9LLN6C+qlcj8
FV388u0c2EsdE8XZmy9uCX0RPmnvMDHc27j7vO5ohLmT5i/u0Jx6pOdWpxJv+FRC
U4VaoO3VilJHoYUkfI/vA3F8A9zQg/rN8jDHG+BpD8Zvlrob5YDJSGD+oGZdRomJ
NNfoKdqDGo590tWzcmY6vYdz6shEj/g5XfWJDr9NrTZ820J5PL5ABo5dFpiz5Lkb
CU2HKoXLq4G/yd/xWAAtE5xOQpWeixcOwM+bhg3xKx4UMRwFEnbcTjDIVFCXD5u4
3g80NjjfYE5T7HQfQhmITffNHns8x3rsqem3Jr0t+DWQmJcSSyFx70AUYu5OWmz7
JE5Kumj+a3UFzVcg2xa/DsNFatVuA7aiJpf+/IadU3zaofxNBN6iQS6x7u5x/YNb
XcT0dNM8QelLaAuMLJhtAcpCVNRFklZn1/wSGCAwJBKA86t+HxjbTG4jk8PUk8+H
BjOuAus3hQewk4wuJHqqNz+g2ukqyK3Xzkw5yG9rz8I9BVVdXBc7uwHOXzTm51GJ
VYbx6WauIF+i6+R9I1i7SPKYDMW0ncvUfIX72MoJDLFZ9K4lUVba+q1clZ+A9BSU
knnFePXcI9CIyHAVkduX2J2O6O1qkwPyIvBL7aXpAEWr72j78BsC+SJEe83j8ILl
Ud+1O6g0RFThz7ngAredGdo72B417UnDUfav4ivxJ4MZ/eVAUxji38on0T2+pQby
SKWihmV8mjDp7HcayDRL1V4RFMdYz8mjZ5PcUZlrZ/LezJF/SgS58w9Ko5oWsfH3
E1Aa9cVL4NtlR6EPuud/X9XjITcShSZqaLQh67YrDytW9tVi1HMsYCw7Y2xAc9gi
mH3yLIABZ4jnUOgPqqpIQb42CR2OKXFfwXjGveIF27MXMXj94lJL0kWAcxACx2Fc
8S0M9AmQyp4nWJrLSjY1ijOwjQg7KOAJ8oPm6YHSjMM4yZVgvl05VfxM8Rj7juSR
G3O6rOxqwVd/I+08ZmDNlPAHliil+hcfeO4S0v2GnO3gCNEror8jomUAGG79ZGQB
I5qaULpruTl9SBUuVugnNTAahuT4M6Bk8DODTu/VA4I7qcjjRCrHOFciDx5k+Ztc
VIqmDExsRLjX9OpfpSBrYVuHWc9sij+RjKP67tn5I/KPrQNvPY/wQChSR6BAu5U1
JA3Qr0zxGMJbSfZAKILVXo2zISFUyqlS2vmBesKRejWWwOXI7U1eFnwDASm7acQ2
bkSAWHSTzarLfAj3cZVl7kPKkKTN42L4m96fe/vQt6J08BUwNQ/agsM4fw2Y3g9i
tdRKTbtKK2uZ50H1OdrOr/Ez7t014nmJSKmRHzRfvlwvJbg1RfZNDZIiBP6clTQY
dlVNGY7YWKj+9NSCmAD67bfBB72HDCHoOSoB2tqdwrCNpTWcf/4AMkNcCtO9/liv
evxeR56RX2jHYEwd5QNEV28+Ny9i4Me1wcfuf6VNE3aSbkS5JzC8gQPOQOD/zkzu
vZWjAqvZpArdfkeM4RFBx8qRbpbG3xB0ViM+KNYVz4nE+NwdesotqPgyCVpJQBAN
lYMjex7Gd4cnP/LZhYsDxLwswym7klQpjCx6Qi7nOy6L/M7zfCjZZ1DKHODP22Ib
b8vNGTzDp8I0ELbssVNGoBR+/a0piaqsjQJC7Zl1sw3whTRNxfqz4mdzfZTY2KTy
u59GuOdVPi1btEBuJKnElFAXH1MWIJiO0+gC8tYWiEwQBNgEyG1J1wzxibyubeo7
Ol6BBHMI7TrLNX2FHbpPib7kOc0gFIM6dVEhhi/348BvOyIFzTvmcbE9GkDr1Q7P
qjPWMfNvxb/AgZMNsMcksVeckn/YoPK1I0mM585oJvMaHQ4ZW9j0vhOS3XaeWJog
gAVLNMeYcRkIAfvLmWO81rc8JZ4//CEKDYd4LEK5xghSDBDXT5B5FYeh4MDCJCML
8gfr+KJvywZlEqA8b9cVKNHsNPKwJrU8vbqeXGxTX4VlFI6Fb2U5kdD/+K7nowds
XIcVYIGKREhFJVFWPxrq6fxZLsi0t+6/fT0wV6yRW3S2YAHSoubYxCWxZSgM/JZy
cR0AyVHQ9Awzt3wSn7RfMNGwFVw0CDxR9pReEpyAfNz+Hgi1OR6LMfX6yTAQO3FB
62oDV6oiNoCXzV8/tMIEk8Shfs6ukHuiHeGaVVs3aFmSjbUSTDs7adNbrmXlYir9
26Cv7HxuSYOvgZPMp4nWPqy5K03DWP3QTqC9vgkRZnwuhGgQpBz3PBhzz3VrDTq0
xpdHx9UTm3xzETTdZo8FlozCdRJTQaPywpcwRddM6FNVsVhqZzQIo8WpKINf0i/2
7juHj4aSXDkgwYZCCuT0bhSkAIpy+yeiTO4cqeyh1Zix8fL2ExBYOzeWqh8BPd6Z
/6jNVs1LymawXNC4MkbaUcP9ecwtJdafj+5+YCqYtOagKziDSmhm0j3fAs8dHJBi
4sikvpBIcjVXvQFh7f/IYDnOI9qYDl6po9fMD4T4EMvwMbUIZJa5E6GdV2tDDNvf
7K4yyPjuKQw84QAp4lJXM4bLM7iPUyh0Au+3xtwDUknk0rezSAI5iX/+rgtP4tyx
G4My5Qkt6/zEowcBfeps3FAosCw+htG0YQjoOjns5smxOSAqm7tBc/c4NQ4zMALN
foT+mUt7zMVbN4qghzbo/xxDl7fEDJCeADJWQnc9pcO5nDlYBrfb841k55dbvSpw
k8Xb2Ejn7m1M7eVszPf2WUcbW5IvpGArLN/hZRT/SET9zmbX+i0wmncDAX03BX9W
IsXSNM0naq4u5Zpk2a577ejzam/aD5T0GALw9AoJhMBAQsUD9IpAQPvD6241zO5r
qQ2eUfBH+obBYBNpHTNH/ThvDZKsc+0BMDqUgq5KTNTFhQClOOg8UNZD8vG2oz5n
aktJPNzWq9cthzrGfrtFe8y0JGLlJQtBAlBvE1Xiej66/61KVKb4QDSOj9pR6ODu
pqgLQzUdKSeF1LTW7/DWbm5jg4DOp9lA3RGXv8GvFD8Tw5f4h6HJ6NBph79/cdYp
TFF8zfeMgv65UdwI3PadZlyyyUDbj/h1JS7HXHdq79Ou9bPzC/9SUR8sfe4hWl64
XbD3qH8f8w0QETNgv55+VoCFqz6rh9tkyTyWtsq30aRsWa+JTw8tiyIU34vV6cr1
7nYmJO5BdFrAfPtNlYHig8tZ9qtVOS70y3SU+gW9YugVzC3RzFp/Xo2Di8ZKS892
qeq6dboVGDuS2qrcBX1e5/mcOPnSjphQTYhR2Z6I82H9vkHOjhXQzsfHn1wVWWcg
Ywc6xA1trJbA5SWs3PvKBEok24Mac+GM2KdQ6p8g2i85rKPfyJ3dVV5M+WcQ+/92
bkMYYEfOryUXQWdbCY+6V4MJkjVIIpwyFETCdwN9PO5BRENoNzxyntB4Bkhm3pre
3W8zMhRvxv/3WsKqTWKZ23EIfhBeAfssDbLttOWXBwixakaFoiOoN2zrCuXIZGCQ
sSlm/Z1/RcPQBlkGtChaTuDJPgNzH/H0jhbkJHiyPztmvzcyNlM/92aPaC0oRnkj
scJH1pVQtg+trFAJfnNi8ZA/r05NUqGRGlAZMngYyMlTmlcMHjUZhfFiHFG6EPeU
4AbVhrSLoIm1dNucxZanQfVH10gokXAu0TwAAHuXFtUb0pMLbGk+oLnR/yBlQTuS
4zyO+TITyaojn9fBNc5v02fnok/aDozontC2Lwokc03POZQzigPqoB3KxPu9fr/n
Zuf4/y9r2AWhintPyW6/8Ibi9yqn4bKdpN2s9ONV0JPVz4es4sjKrbyuIo0pqkle
cXMqZRPpNdZw0X0UiBrY753g+chpn2c/LspXs9Vxq4c52bvBCf6PFLEoH4yfzEZK
H1PFItRU3PlLs+7FaUL8PPA29z9z3EkclcObzaaODiZ1xp0BWwYB+PlpaTpsT27B
iwaVcqdNjCjxrAooaK40MDMY856zNhqbkNAuf4m8CFiJPeQAsttGD8ItszCC9iZm
2Udd88alrhO8rITGfL0UZgtXnPshHgorEE+dqCUPQKIuF6PvIw5hYxcV4Z4RjePK
kAJMU/jxrBzDcgOBgyIE7PaNaCdP1rKleBSqN+pZUD+NXBbscx2B0C6paQamgUvs
yvg98jq4gJxg3KEeNZGhPAdi80VdBnrjwgLVPQ9fS4BaRm/B58fXfJGqFoM522tM
dN49wRFPyHIhTZ1c5/gK3iEtxhWImbbNnJrnxs/2lBjD4syQkZ66+8UFO1K3sgBR
PkdIbAZdWQNCI3khGAPB68kHLpXIO/OSIXesBg/yz1VgDPecvExwGMzdupf39LcY
Tt3xRP4SnEXA8ekKITWaFMYURVmIgxrO4ehJd7+woPDfAw75kbkt6RjdMzO/StmV
ykIDfuJKJXSNhPNV2WBx598CJFnphWY3tktwXdBgqpi36Kgc9jlX0L26cHB7Hcv5
1QP/AUMKWrLTvFvEL/QYWme1SZcwkZTI2NOBE4HikQTde3Mt6KKjr6dzz+N7q3RY
DyzNXiQPTTRd2sL64IsAmZkI5ddj18UHpuvr8H36KoYZR9HQb4dkaXqeUqWRYOX4
E3MysHfHYsmj5Vy0Qk6XDrjvtpkQ2dChuf07T5rLfSinaPTFbvoqt2hqy9KMgeWL
uzLDiAiliXwTY8IYjk0R0B9xgupzuxJGtzVeRm/ENehGQTYuVtm4MQAhNs79pPMK
MV5pPiBeDCN28sYDrJJlvcwCZAaYLrK5EDPoSfQHZhKgn1OJ5msi4YxDZEiBuRNd
vyyo/9Yir4TRcGwIAjsCS5cKB6jQp1eql/O2zwEmTo47IY9c+I8fNGCvVmFZrYjl
1wyyyKNk1NjCtoZURRIhWeMKeVhgwGCn+CKAp6KMC8BFuPJcT1e56czlH/35ygmE
WIuORXEXU5xgfQrb790hSaUCDw72f0ifzSGTZCbMbSvQicsVWoyifmE2oxuHU44W
PPEs8i8JnnwHcjdEv/JCZUl696zaO45Csfgj8+PfXCnNw+B1gblaNGKInsCaujvj
sq7VLpy0nI9flmv+auLoegNfaHWq0fzj5T1zuDRlPAkG8iIDvJXgHWAP01uWJSLb
sC0t+pcdA7NUNHRnT7zbJBmPmvfd8Dk107RGhCuVjCAQr/txLoNbx3+vVDmY982Z
zVAD4xeglPfC2zBMvETUN/ujkiZNYL8U4/Bmn7IrvV9YqTN6O2679FWqyV0aV4DX
yqOt4VOoZY7fuUh8H2NHiWPBqOwrlw3Q0HLHnLpik6Qu1WyXSpAGdpNXDWoWwzHq
xwYxn9YOuHXiGNP5N5Ro3x82jD4jYOYrNaeWs43NrkDOAYA8eM4mJZntHiWkFgZP
vI/QrUoU/mZ3OJtCLwTXYh1jpB9Vt0TDjNqKAqmCvakbbTOb3S3vQOXq0licAd0U
82XcFyB4E5IHA3Y63LuR45CbeeXh7IVwM6DtHqt8CFlpfw21DWrdcynArCiMjQCj
WMfgRdp/qaykYUxH0MXO3teDkv8CUlUqlYWJxKmEwNoKJA+ET3sBypJtQd9AlN//
XnSGzU2HLBctIwh3rjL3O2WjD8i3GUEEX6GTJRnb75WLM4u4JAUYdRzfalP9BYlF
CQen7hx+qVm0ivpF1lBqrQRL1tSkhqbhIpipL5yzzwTSqxnQVUYvc8FIVQkmMYWY
gmvrjJgdYQynjfLBWmOe/PFB2C4SGdU0d1hdO8TFpvCMKUpOIcfKdOiRUkx35QbK
/6YCLDUlZ8eHynyDVfo0hRLYn1+T3fNFeuwEwKHyYAq/r6efHMb78IALMr17CE2i
8RFqodyibr0ixZzpf0an4cSAKJRHXWGm866mcwMTaQgT0RSaA8xM3CocZSq2sobM
qJ/12tvOZAsLxJ4VXJijikcOH5bk3646tskh9kGjATD3yz486DAcHOpBLn0mRLQC
c0YJAf5+SoPCtUBc/Xo6gucFF7dVjnisIMkzuBRwcTaEV7VqLcKnw7QWXc0IyBzv
bonqoSqOHgRHHyMYcU0V2ZB1w4URCe2kX3rqpaPev7mCGL680mPXDtXYP4hgG44O
O4sIVAbMeBhrtFJUnCiJMCKV4pGG0J6vAPjqpWuPk7lX6KcYdKaPyYuJX1YbmJd1
aRmbEDLoXfC6KidpYPK98KD1YXdwsLr2HlllQxiK9q8Vum4Nw5UUK4QH8Uyragyo
mTpvC/gsjmufekUKDR9E+H0hU9lP2O7LBZUbvLeKHkwqeuIdDhwJXvCJCpR6seCz
Z5HOj80IrSkbn3M38vtBDjjrK79cOj7SBwHJs48hZynnwSW8YWRDHSq6nhxhzW25
JB9yiKdv5PQ+UTstiJXZ4rJuD8ykDid23JWmgZn16/6hFDKEehMHWWc07esKO/tt
0B8PeRVRIdHsVC4LOPP3v4WcdcqkWiXVRnVcr1ARJXsWQuS3R9kc0XaeOf+t/cRi
tKRyVVovxEQdJysrvDPc7oiXvzOzBOn6RmaOr9kRFpScvRKwO+VQxmmYSK26Ysq+
m8tFB1JiMeIRjH1tkoFHUurIotVIia/xPJvH4x89bPZ49DV9pBFjKnDN5fBJghw5
K6QehSPB9KR0xVDdlvfC5IjgTaSLQda9qlnUcArTeFudDftAQOsk8apxkA8i86sd
AD+xFNqz7Dr6OHp+Jpi5/i6s2giFUNLDkx6WaaQoc/RNLQjCUUcEivwM66tEGsXg
NsUno6ibW+YnkjY1sEgx/AFe/2GkYGOmoiqH6ECNsCqHI63YULa0sFZLMep6wUJg
cFLRjvpNx0XeX95jpTrKzbYlICbI0Jq0ZJXBDAwB7QElpSuS9nyOe0izPOzvLjt1
aAV2VmX4wdHUL4BWkQNjj2OfYeo74bN5v7QBhwfyRVfLcRc3SkvFmz+0ggfsQSo6
ndagauKeDqYPqIAI29kp0rkKF7eOt2g2FgT6DFhz9t6b7L7qpKLC/58HUdfiZFB3
unw4GSJV9TuIJuJ9lirBAP5AfqdRXvvUrbEkD2krk4xnsm8nIF8qTwzQIHhcyVG2
AqAjhYO3zgYx6E7ssrXL9JcEfNe9C/McdAyTtem2wO6se4+OFBH2VZNWSP6tTF1q
wC8qXMbRYI7Daovno1de12wZ1EwIb4MYq7AqjS4pAl78TxMclF6F2fqcBaJShPWh
vPdIJ4Ve6WWu8j5nDGpEdl8j+VYOMLcJTiU9bd7oiLRKhzeB/tVAl4kdUehB1PDi
jf8Ki46gvNR8gBZAPew31VMHYlukiN/3/iDKTUmy55qTFL98rW4TlwthgevfnG9p
N0OSpttFH62Haq4PbM6/bfrEBu4hnvKNqEBW585tMYLlTBMEMxdb21ydQDhhig4Z
GIklzleKnjE6R7T2NQQqiXQfH82sbrO5QssPmWAppc/YykvoEyAoM+ZkBKvnAhNl
asS/QR1Ge3ZU5bHmZnoEIKAw4BpDZ+WAjYYAz5CFFC8702Cz7+6KUEK6J4FV208I
hvTXyf5Yt/+DtRv5XPnKnubnDkaq6gtEP6clqsJKf5gFU8DtFOjHxn6SkACQ0AGp
jGZHuk9S0jYunvz1IeVmPDCLtWbSWEJKhpphrMuuG8I/1aOwda7OK2EyS69Q6RJ1
yNB8pGGrov0x8q+speKCi5dIXWkZ7V521ysE+p64J60oNlQZ2dt2KOo/9YkW65xc
8eFEHBPr1uyVHlLEzB0WkXx0+hV71MSkVntg7j5xS22QobDuBeVB7tdNig7Isp1Q
qrEAotisOhSjpNHa6i9CQgiWua4bVAwhVrKdFs8fx9MPixZhqvJmcnGYScogWHME
pSnjJEM0ygFtT5KuE5nYO0rJ7d6tM+2QIIkUmYirtoU8m6GvcXHSBDKO707KHuho
MTBAmAX518ySO3O18gSUNe6CinjDOB/5jCdEykkxGANOV6dR/ZI08lVTEkrESSdR
CvgdvlHuocwV0tSTv1agvIh6WD4Boq+QgiQSzGiaUSYviqjQRGQmZpeMBKXGYDE8
TgovGFUtANGH0Y/FVvmpeZ3ZW5PNnusjsas/3guPdb2isFpNFEieV5wdcGOrRtUH
VpthkLF/UNu8gFYY/xhqQ3uN8S46yPORR5QWaP2Sff3D4wvch9fzqOiEcX1RWzO1
r0h+kc23iN/1YurONk8etCbIRQL3Tft2FZWj5Fb+ej5xK6nEsZJPwEkpjarJkrif
CCrDs5uCbPSXu6DAH+/O+KqmloWW1HK80121Nw9BwhNEF7n1xh1RHqjsHdOF5FBt
NfoWh5/g8VSCKsg5onZi5CS0xHfxj2SSY2IuLlmycU7Ws0yPXJOQkDIR6fKYFcKy
szyhuazwB+QkqaGIOxMQ4w4a56NSK+3YXpHOxBtFC/oc0ndEYK29qBVLZ3crUB3b
i86XyC2jJe2I10EBNnS+7sS7oKVuyupXTwTorljuaFCxiggEN8+ySXt1jjRuz7Ps
5rBjZSHwriJyvh+yUITXpwT3NpJ27jz2xVh4ETffGp2Wcwgpw8FszkkYVah4BtHA
pJe4HEdihGN4Q+27ii6a/nuE81GGbJwKd3sIvRyz+lH4VrPKqW4ApundT2vqZEEY
pA1gbFZeLOBDo3sQmEKYf++inGbmTdcaWIkcgplo2XXQn1X+bFF/EtGPg4GzqtZE
VfiNGqW6+USunNtVvVIHU5IgSEbPOIXCgXCObSP97J04Yq49v2jSp0O2UTOJoXXZ
DfNpXnu50Wn34BAXF4K1xsBXER2rGQB+E7gGM89efxaH48onmz6zRNWCLNLPB5+9
GYiO/NFDf0Xbgj5o2Huqsz7sMnkqPMfJUAuf0LqcX+KP6DS0c2ZOtphVvOePqH/6
yL/J5P6hjRyIQK9aEPFV/VBUmT4E9otV7NIvnAfL6pv44JaavMWT/ghbPhTpoT8A
ugx4vzQJnoBEzbXMLkQPXmWhHGfyoRoWMO/64W7v4NQoMHYOYZ2OJB8PiV/+yaaL
p84upH0/K/E81NBqSwGTLkNZouxt4mkVOL8qLZvr6YkqHF5taSZQ8fGmrtMGLkif
M3chWWJkpBlarS8F49TcopMTihzOPnR/hd5+/yj0ZQOEobPs2BfbGAG8o5Es0Lyp
loscx5GlXeKAJyGrWD6Fvq10XQthw6FSec91bgV11k9VrXu0iIOkqIxcoZk+WLFh
1DCqPPEN2NsRKP9XoW6M05qreTKyaNDc+V0/uhB2UQPZhJV3NwtDAXVa9d41ynMW
eMiQyWLpbLEcYLhtNiyEHYSqrf8XbpJeBV2RPNI6JCzjGmffVrCYUDfYIDb2oVX9
w9+zpb8r7oXy9AU4JSQTYvG4ZT2WpB/l+QinTKZTQUacEtaSLbrLQiuozhzsuhfR
wnz90w3lgsRGkFHmC44rLdwW4XqiRNGcfio6TD6ox3a6mHC3vCHG5c3G9zWYHraN
1I3rnSUtvrQq3v9rdQ9NGbdmpP9xYDZIfZpchhXqtIhgRYgGcAqqe5tXpTY6ztT4
JeJ7kCl/LCOiiEP6T6z9p+6A1QFxeij9mcQHyQkhstlVXz0SZ35Go+s4KpaZjYoY
ND+HvX2XMMYhFgjdxlzst0tklM/9zHI/X6WiqPdGme2ghdaPuJzOzdWpKoTH5aXF
0IXng425Vlji111husF+oe5UVYZSTOnP9dVB34fuxHnNY0SYolCeyjQBzTgJTSoF
CRmmPzncbrTgM6mkGHj/uKtmsoJkfebSd7CkA3h5hov6yR3P4W92D2teEokOFPVi
iPtZHXNPNr7/Pnkd1WDD7QN4X99bTn2OVmozJ2BF9+P1ppymR7jq2C1W+Dt31Rq2
KTfgo4QHoc9LwCRd1W2Pup/GPwpnAhEKM15BeUSpRhavoUYYZQCrAi61sVU91IVc
bEuPRixOa3KwsAzFMA8AM7xuUyu6uBJ2mf/FKrmnodhBWLHzzJShkkvVGr1cdHbU
IGMpocxUybGCtFCPCHy1DatRKgLMNkIpiEw929GjW56LoIdyTHDyvylDfzM/Tcc+
kyQFLbm30zszTqdEUaVhgmaolWxBJVstAE6y3csuBrFQMd//EqJd31bZ8XIzNQOR
5XpgTD7jxhD/0RQaJ/D0k1hdeUTwsf2C9KGDCQYrTJV67qqujFeRBmtmHy0AJS8C
PGhc+9jPS33Pl6sumo2DXwPYARyvSEr39DYVkZvgxHXbg/eciCwrlL5D4OGF7TI3
vOeRmqe/5YqmzVvABhU6hgivjLpq5fei661To3wYtdMblzoSO8nmeyH/vAjHCjEQ
uZyK6xO1QmbjnskyLeiHerzijTKyMriVCkZcK4sGoqr6tPkchMYrJIkPLN+f7fPs
ettKCd3HUFjLv1o2p3YrzyxKl+OjjAZ3dSEnwEkWT1iABCwqwavv9DMWbH42Q814
29XqSHBtPSWL293j//R5Vsf58uLgvWh5KS2dqERYlELaazHLuEQ2pBOxq72ovPfS
JXmPsYQPlIEkAm97qboq68OoB1QQiqI+0NZwDFEMxImfQIsD7jiv0PqCNVFNXzCh
PplVK7WeqHr4ZhM7LvAfRWCDHrN9jk3bbrqQS0xn4CNO1/9q3yUPq+5v1hmm4RfQ
3DVCAO5sN4yNhbInqqHWQClcMoaY/IQLyvdqTRhdFDHDOFo5OQxi3Zy/LVomYjNU
32dHHSs0iiomxRzJFO1lE/SP6fQvzp85opmNhBOR9RIBgshgKO8hrbvlG6U/k3HU
CgDKvcuZqRUljJE/dDRBptiqGOMj+Z6tJ7HP3qMhTrIGG3BEpzmqlaUICV7U/DiT
9RNCsnFMvmeAi6d7uBiNAxDq2jglIrjV7BAGRYRUqKVbwNfHQ/uoBrNg3TMcAaLN
NCk0YrX7wimHgStWz30zb/mAl4BaKE/+dIEaVn2HYdeo24LtKTvVPoFE8/uJnAHP
xiFrrBLZbVlJZ+7wgBuT6UufWMQIUvhRYsfLDwS5dUUw7tTvDYgTLwtUZ0zTd0B4
yUVwG17rlyIHXhUFmNt6eyIm2V6jFouooimJ4Ws2AmhSG71ut/fY0bToc8i3dhy+
q3qYcxsda5HOMmxTeeHgTlBAf2OBIpmoMx6u0WIEo/lRXK3EagT52NWicQk4KPnp
bUjoJltWn+6O5kolnjJ2Y9OSVN+QYMdk11xcEOV5fxYx+UDJegdKeMh1vqVQ7nnx
hn+7qy+81qAU+X5jWQOpFtFr9gXZLyV6vTwBxA/yobbVmEo4q29NXnGazQ8oej9C
EiKybtkmSxhWosUkRn7nJxxHNBEJnc6LTkarBN3efxU/eNT3BjzW2XGCZ1Tpp+dG
nemkj5p6d5I6Ft56YzIUEjmf92F48QaypYdzitI1rAhHJ3OSDsQQT+K+jSBev17m
EeTwbsYfnKmW6WuOx8jvJJyVT7/KuiBzILGDUnvobG1wNR3049XO6lQA5wuuuy/Z
9oSmByyU0coDl/n5T2o6/XMW6AT9rithZ33ReRtYtKHK2x6hCkXSFJ8o9bIedJS2
K5oQKWvUIfvNNYFVTC9mSeZgo34lWwE9sNnk9VI1s2mCTUSIA2B+ygsF2Xz8o0+K
zpFzM4g5604MT2AnDVJH8M6xxANuFLWnKUNAqN++MjN0xqFzJ/RpkrQDxKx/F3ek
pMz25ySvhYprGYzcqwJlamk5NqopfLqvAUTUkbZVLuTJ7HOs86umKy88sSXFwMQ3
5WpCQnkNd3M7pMygkD56DNAledoJookZoMJYgLIkq+Jwn2wnEtM/WO1YvBAagsfm
SqMpJcJzSgMlA+yJitvOzzDxwiqLHd+Wxz7Oe2j+L9B1eF0znUHeTr4olxx4YJyW
R7K32FAWDo1tjpA5X+J1fmA57vAUBERPM09nvZ9YhNXxEHTXc5P89a6sVRhZR7iQ
iL+r2kqnkziXUWb6AZTRVQUwhjkHxbL0sqIEAbckc8UUI65mfeK/+GbFn3taHOIU
qm6WHU8Nx91MZmrbOtlTn5p4VQRLaWjikhcPLfgeNSgbEKx9tiLdZ7XBBaO3t5JN
bGOtAIPP6mZnv/qAjG49GgB1ezOIlPT/q8iN+496FUZyt4zuDwMID3MkX8DLb4ld
1ua2Q2wiY/pWXxvk+vj8b36ur6sgAdqblzln68V+a4w6Bft1VJEcipcJ+I3T/jMn
EBoZgOvNo9Azwtqim1maocUh7qezN+sqYhTl1jLWcIpFYo9TwbCi+sF5bNssCsA2
WMtx2+QNpF2yvnqtr87SeR6d5xL/1Vk1+iX1hM/swd1M3Ki7jN0T/4k0w+ujNuId
cGWfNfevFVluiZqIef+04DLz7+uP3gx1y2AAfUxyuO+9hO7HQpu5+u4XqwWgbn0U
7CxSXVVPTekXZNX5/C+CqCmtlGKDFPs64O6aaI4nc6e59Og6WvQzCaHFaSNGM87U
2hXCzEpjSlJK7yL0SL4vrUQh+xxpVJa6hgVETVbRyexQKOZr22BSqrdWORMHGfyU
cXtSsQJpWVxQO56OkCwNTdKJNUPKFdX+uBKiR2fZDpBJN+zODjBQtfPnIeQ9OkZU
BwS/E3MEUAeq4Ln59mQadscuSEMAlpw4FuPPJyn4Yuuj9l6en/jOVZFVeZn5GVX3
4GXCsMGrKwAq2zib2g+ueLgiBingl+4d6zFepiunEQrSFCHhZNNaWad8fuiW/Iyb
1O/2HEGYgFoaWK25l6mufAW0xiKg4WySWSEPlRFuv4SZpAn6bj8DhIamsT2jjp+c
Ts7a/kY2pVxMcS12Zly5BsDpghSH0qrnfA23R/DRZCpCyqu1A11OyZkvKPvOE+k8
KIxytbYhlSmHJhnehVQENfCllqsNARJO+p8Oug5m8faJvTOWk86CfWFz2psYHcR8
YGAO031dtJcJsIy4s39TheKOuCXgxZqvhIX2346SEVlLjq2x/FXUfkGPMrRHUr9h
nCbWuiSEujk/axhSjcCHf0rYs8ZaOo/omCX3QnIBPnLIg9L2sevkUwf7IgRFNHKt
ZC136EHoHMWvR2iW2twLyDYfxEZkwE7Ucf7mz7aLU2aryIhoyh65vOyZXn5o6PbM
sNJ3zWnp7FmkblqvYdhX9KFzFhAKBDy6yFXQwkCfrjdfCMmFFnC4fMD+rP6EankM
cOgR7acziI9AOCIEYxmH9V6bwfeYKUx9HrPKVBou8BF0wEXgrkt3kaV7hvR9BYAs
K1hUbNEpH3qz+IVyUzWdVQqeR7fgtYQZvctrSEyBF2lM2ZXLC5gDduAjxwanT+uP
x9eMRIRefuxmrVXTGS8mZEXnlXuk2PGIPXX9oM1NkAw7jgzbM7ieUufy8NEETR4Q
BytmohBr3pfEP+vqZvz7/D+70Y61NtX5xwuRGiSPzltGht0Jm3noRID0YKMM1oqp
9WxVTW85JN72d9RH0PbdPzuRbVXqVCw35lpqvoFjx93qAFOdkZRaG+Cyw/O9OcRr
eP0ArXbhHdAJnJo7N70hDxtr7ppbi2X64tyCCnkuCtbCaQlZk3HpgJoH62sRtHWy
J3mABA0LQn3RG9AIrdL2adzlZBHBhLpeZvvRKo5uLRIeDSWbDXHbJGlOqU+8QUlp
6ryq7Pn0tsp3gQNkiu09U866IwCVSIywHbEOrt1KNVjlWEhLiXHcdqyNrV3uBlMa
m7b2rBBjT9FR0RoxAGp+LnXRZueOGhEVmBjXO45ReehVg10gj5txEtKHq73SKZKl
7H5r287epuKWaRAJ42obpmKxY2JUFPm+p8wh6YA9eRtHWtzN30zxFkJ523TF39/9
0kaRE1MNDhpr2TfjpwPKNfw+390GZvYibYiihLlxdYrEw2hhvQ/TblwqsjA3R6Mp
LGbx4D9+eIvDoWS8IbYgOhNzQWAIjMz01W64c6So0kiv6hHZLktNktyD5X0Adg3b
UF8LzTtOe37mE9hwF6fgBVT038ZJVDZiqGJ51IQ0lFqsPkmZ3zID5Pm5TT2he7Y8
yFjODNNHHwgmBLA6UrDFc66YXoPdFieks9pGcUFlK4uyAwHeH92+QVjZOCntgb9A
/egULeeIzuP8q1Zxc/UAn+5tlD5SGQ9O3EOcmDvfohyTnsLPaapy5TSnV2iC5E1g
+RpPE+925gC6Icw9YjmpKr9Adj807g6eD3QbrMdU6gfRlaMfwxnS9204F+lL4nVC
xyXMXxmn5scHQGKwEfznhf9SkUF+/CdiipsaGfApNMDWx5N9IqUgaYle1IWykv2b
072CYxM1nqMHHKXHu9Tm+fsYqvgJaeNM0wA6etbD3gJURkFznchYuxLiFT5TKXCk
29chTEu2/gPgm4jw1mLGVAd4VZz4ohC0RybdhXwvpixhtdo0aCR6d9wsrEfzlute
WPsBOI/UYjw90q8eP7u37kpF1AfqQ1+jG3rqq1CsvUit5T6ER/HM/KRHTh6CFyAd
zRbCxQYzjDYkHU4UPBZ499RLRKr3MWy90Zpl6+6Z6w5ERQOvle1xRiyaRHo0Gllg
gvMKP417X+kjytOkX3AZplDAbL2OFdsx1hIaoVkMVM4Du7UIgYU7D+aGM5sxpV5x
yes3CYmY1oFzfn9azQme0OXmOihT0EML86UAYRN3dehP5jxSn0J6RK64TMu8QQtS
/Igsj+ehC7YGt98MGdSsOADC4E/HbZ4oEIQWdl4MLMcDUHVK6IQypEdo3ZtQ9XTg
obrdNb1yVIWqm5B4HwruTbDcs73QJMCY8hkKCufOtKGM95LdTWimi2KFXL0j0YHf
JXU2uim6evldkTlLZP16Jdzi7VbhhbOzP2/xZup88QstA5sxdDFnBTLN1m+4JMNl
UrXfP2I9Dlg/fNQ8Ajo0QlfDCAx8dn9WzST2KhVVZCYdJ+iZ6q0qB5GPnQ+MOB4M
8s6or2cTP7BILkLWLSC+fQNCf8WWzWiVR8A96srS5GoWuG0uHdCgyFzLsSLPyqP3
qoHYMmw36bbRxj1yqWwzp0MD2Q+JqFmFbcnEMcsxKy2RDTM+hQTS6/JW9rESDRq9
UMsS0DJ/U8ytVI5hKd6rb3VCgo7ONUIgs32gXhMNvT0nR0byLN/urADdq9f9kW1S
rc3Oqe54S/OTTCQRZJUswJ7vtDeSAcw7Ttvj06xdBCFtyTjeFn0JpFBitjz/4Cf1
vOZ754gcxYZi3vxmN+tPS2HwH+DMVhbabil8+buG/kO8WRiAQBHowzQ9Xf1aGNFl
eW6KfK73FzlvxsMusE6RHfQjOzMpDei5i8G4hQ/HwQM+TmlMgH9HmKr34sQHppDJ
kjtJYmjw8DFP4vcMwT6+Q2aL7LGvKXh9Jz9M/J9CLSFafVWrm0UklJBVKFy2b8Po
kA8y+NNI74WA7OxE9KmbelTKbfAloD+VUOygi2a/ZvJSnXljeWI4TkxG4lAPNgSn
ABtc01Xd9kL9p+Abf/w0wkkli8RIIriPfy0EU5BwbISTaOsgVwULBa2MSwgpO6Ct
ufUCMzsOO4tVLMEbgtl8itn1R8ZvMu95OiFyWwZXJNhzc+a6SF/7dfuXRYspdv95
wlNzhf96U/va6/ec+CYsVa9m4ywliQpL81AhfohzWfXNJYUZ2ZIQtcwtKwyPNCZG
CpmScNeLvcIKST/VDZkY7Uvd+pDF8gm3PUU6gGoBS6aoS0joSDfNUvbdOaQUB4iK
ExI4zEmsNBUhPIodrQoz2aO74WLlopUUWBbmPM49iJsi02TnaTOwrS/EJY0NKdWy
D2b7kWsp0Q2WE/ZNtE9vlSled+adUXCm5rAC2t8N04+JKgHSl+v4jNdldC3DYlYq
rRyMnjqHqvzilVPfyxsIz57+fbZnXboXRut2NRgFSR6/HqWPdS10+WeMEIk9QfuO
AW++JMSaGwhPuEsW0Ri1j0Ekkt4AVDdZsYl4MUDCa+zREQPvnv8lHhnDEN969+OB
ldRnlgquSctHY44BJ5vcEG2/dGD08sCrWNLW9e1qclvkjviThzL4NquE29ddh5tI
mFLJtj8rFTG7jw6tpazAU2fibheK109JGwD+vwBmsfHmkjbfDS/H6osVpP7Gkdzg
oA/+pvtmgFeDsZlvKSFyWrFfz/I7tntLlpyIHuoV4Gv9isG7VTMK1Z2/1aHFlnj1
Etu+PtzJiDwMJlDmiz/NZ0XwV/eHgdMSZE1p452FeXyRIboWDA2IY27mc+RasIRy
V0Z1/Bm4anQYPqyNnnmRalzTqfJ6VO5r6p7W3hPxKZS2GB4+zTAXRhl/9IIpDqqj
SAUcDoCIwJdX8RqWwhGZzHYTMSXrE7XM3piSauI9vY2CBSeQLi99ZxvBbE6L52qx
kXq2p+2yV6QuNd2+xfpctJrs7v0n8n3N54ZeG12o/bkbRXwqqpfSl2ByGogyiPgS
2/fre3vql4QZfUNVlKg3wS5xvaKaoxcaq08Ja1yFWHEtsY9BAMJQFoUe37qTEPFQ
/PLzUxGs8C8rOVJuL1DMCGG791cc6JrMhHYVM99OdKCUZ/KQ0uLI/Aez+vZH7s9p
9OeWrKKUlX99aak3yMOJWJ9qKzZcoHrxdGUZgjWoF+3ikZ+m/lAQg4JZdeO9SKw7
/Fg/sjCrygH1MgY5fteZwKUDTzA+B0Ak1dl3KfbIKqVkhSHe49J/kpe5mJhc2aRS
mWCbyJawqT3/PZSViUs5EciCwKXKaOew9wkuOJE393Tx78jDqV09dKAQtXhGv6Nd
LvU4m7tOLBebvqTEMd89b3Kk9N8A2ZXM+uYjI2rXdDWZ5whnujEoMJK212AqWGwj
ztG4n25aYDOdhRaEcJwHJnbfoCJc8qOgZknqD/Xx9yMFH+Dmt2Gel8EvcSxaCgtB
d3Uy4xxMpKF7MaJq7LjZxk70Iidc16gocmttF+bpPmBSfCcTAqdeIz/80Xnbmqi8
90O6ApUWCyYxr2Fh2sAvXK19/fVanuy0UX1zGMTQXGC6pLf+510zPxWAu3leGL1b
XkANe8L8M2b0KCqQqU0qF+5sZzzeB1u4/a/vwkcZywa3sKx6yjG5LTDzvIOsEPNJ
5aYXDtFoTyqKOPT7oflqZCSPOJ0ip/6nq0k2PEaizCRZYmi3n88TA9t8COPmCUva
vsLuHcH1DR+Z5uECkxsqfCIrq9vkP9MK4RdbXUwakfgpSztmkKjKBjLcaiENOURk
yVK4TGQTeUs/BVniWUL7xGJ0VHcAi+SEI+PlAmwLggkxTJNSliYVvO/As6gj57Of
pkQ+UaZNvBilkFe1jlBGiMIWgZwu0ZMcg+XOnVfKVk7jRJWzfi2XTO5pqYFf/J2L
j5VIvvQMyEqHimyZX5AbLgk53NQ5bM9LsORiW9Rv6hMmzausK0jb4sFBYPL3Wley
aOUTAGKND+nuaCntD8sDu2P08jeufm4xd2HZDubiCTLwFSy2Qtk0HNiEcfJkoHrz
pTnAwqSgmhvnlGNosSBXr/EPEoQIsxr5WRaeCYkrJTff0t+1cKXITr51Q5+Lv7Az
EWFtCUUUzwCw0Q5iw+ATrQnLCdTkMAItVQoiHxavncAUHyoOEbZ/P1Gq11Qd4SwN
6dlXNAVSoaNBTefb899FgaSEBRsQuUvygL5YZksO9uLbIIbEY94nHk0z2Ntmc2vp
JU+m4kf3FqHuDdotc9uXUUiAncqMhpH7IpdNvyYtLp/lR3BWMWbI1VR3jkyi1fKh
TvQW0YzO1hM9thp8Eg5oYEi8W9N8ZT0pwh5zXdp+LNWgdQ7Mx+g/BrgM/PkfxhJZ
WFurLfhDnuwbsHzB/FEHXE4u72QpMX8JJO5wFHVQH45diybs48MTHaVLSg0WgLNF
z6m+LFgfWFUGb+unWsGDo1/gPMRzq8dNZWg4CCVZQGjVtdT7mjriG2CxxxeCZBac
FHedJdUlBcpasvXGDq7oX/YdXgPfqH2+E0ClWZdlo8rmnrXA2HW6Ls/VHcwKX96V
UmZfsxmqno/+01c32lAdWwWk5tsNeW31nNdSLDvUPAsUq8n5sNsdycZle6ovFDqv
07NIq9PBMeqeIFOE6tgtPs8hTn78MdZSwVE7usbgbE3UNx+4M15JQiiv0K7hyqan
/JdEpmNQPPgSCKqojRoxqQlxrlPUUJK4kxe12QzdVYkBpcWtoQLevqpLsUhP7hZE
T9QFhM2ZwePtg2EQ1+AT3JphTvVNogTqBXjAUaH1332JdmjP+vevya8MSVFdPHDk
En5bo9vuDH9BaLOvglgHtEmPo/DQLQB5GYlY8uCTsHyDPsKiGhknZfvSsChiKeq1
5OEzP1+TKJ4cHID52cb0FsUdlMISNcq11PSFgU/KaSssZ7m8sJwVzqpO7YPr7UOM
K+Q1OUpPewq2gKw0ytaIrImzvmecYC2GrXti9jWhStEBJoYV3kHOfspHzeoTeZc+
jgoDPx9m84HxAfeLVf0DIMqMlpa/Kxom+/ZtAWwTitEB6PF0ZDssYAy/WMeXaRie
Elena+BPzDwOWyy6q0e2VaDrDsSbac3OC+8ltuoAf4jrD9+bCbUYKcDUclW4H9UM
aATCBsvhgTnxZjpTOdAvEI90oii1inEXU6NHjMNkT33df8XbznVWKCga/2t7aGrr
fNWQA3THQ7oza4ogOTbJjJ2nzeK1m02UfovL30bMp4zNvr8sm6ja8pVvyB6ckOPz
n2HgY82W3MncJdBf4HQ968FXIvqmHzjfQzrJdvoJwBIePF3gYrB1CEuxZUeMYiAT
BVqHL4uU3BxEw5FtxuR+k1uBGr64rY/Q0jki4QVICKDzQoMHmPZH+BtAVy690fR9
88smn3ZxZbgKyVwo4APKCAt9Qqh4zBBaaEy7jv0/m0WdWKcbEZsSVTxZMpUh7+TH
BdjH45d1ZDk/0YuQ1ssKTrnDVBBFPKVz89xOdrqSSwQVMn/Ae/c4OQantJCnLPGX
oaJezdLXnftMj49tDOxV9c5HQFfwUHrQqbFLK8xoPUqzbrbkGqb2kLt7A9Qkv7Uq
eMDZeSzLZ+v64FTijeEM+QNLcpqKeivMoO7swU+FgRs5a9vem9oFl1hKr7KNScE1
AhfienfRUfWs5Hazm2D37NPkVvmLx0rDNroOZnK86EFBHdICIQ73ooO5r63KopiE
mLO1zaSCpWvfdx38SnovPpXhxisy+h0pL5PSEjjEVjrUlJVOI/fIls5SK3E/LWet
rsnQbcevvz3slByEMEiOX4Ae5eOHRAMrS/tVyjiSS6b+1j/5+1/XX+4l0No39WHS
DWzEVNgtFn/Wg4jJGf2XWsG7Rn1R258/kVh8A/LUuvc5i+hhEXxHxvRf3h9Fk9aK
DCqu0BuC70cJWeCoKvPSM9c+yOHiZRzJhfE2YirRv0Y0hJj/HDfzpDCPZUxpoGWc
rfj7KVdyvoB1QHp6c9dOj/VAFpQvg5DHDJ3B9F4TeuYSSqr3tm4LAa6K3i5gUgr1
D3bkTRKjN8El/CD1oNh3/W7EY28rFhhsGorwofTVGUzxMo5TQoDBF/wOuJ+neMoy
wSey2vihTERWcrsZg5FUSZ6fTCdJnlF8logtH0UbTNSXRIKySQM51MBQdM3BdzvD
kCEj1JNzIL+g5awrzcoLCELIMmFgXcgVIzPnRW0kSnqn/xS6j+98/EjyYutfPqxb
SbfzOCaJq0LnEdYEZ8YDMiqjva5EadQHZJ2LJ0/+krNGuqrmbe6bGW/BnRJT9n9/
i+94wRTbIOnrHAAPv4a6JXJhVQEE7vBtCVoAP+ZJ8aEpyo1llQGlALYgL6xyG9LN
9Hg9kwUn2Jacf0cxAJekfrvoCNU3yl7pu+aqsMhTonDekLCTifeU/iH2LtormyNx
w9OXvI3sMVql44Dz7Wo5YwWKSSWPsAhCTaOwhsqwVjr4qa6ytWEf/9mxzLEoTWVR
2jrSjCUyIZ5BDQQ+CeIiJZywlr5x5OzSDGywegrXncGKb+n0wDs/e0dSOwfqKZ5s
8cB9Td1LXVwksRuaWP2NDU7FBxoihS+di5UnIZnQjRPcwjlZpKCQIeWKEkdiCLts
/NbAX40+J8k3XZuqXMQp6nHHUClyYiKFRpOskU6TjpSSP4ExGfdEpxA+8vnws/aE
gjLV4NjS2Fl3KcJ5xywoBy0f9Q6adb7HPU9zqfnNa4mBEm1SxdhGSoN0Q41ocwt8
cr8tdTzFNtDlIi5BjsUruimU6W0e6W5DeGJfu8u3XLAO4elor4Vw/0tK85AP8s10
7a9WBYevP46YW/aDjsiGm77tsULqJ9mgdP/t7XHM9k3CmVrw8bnE/zVEI8Eyxv2l
V6/q5mEqse2JkmVugBj2W8Ja1KuGMS2bghhd0LPeWoxF4Exj6jeA1IWqorx/922P
yeGhiIstxBgFuTrarhFYxrhEX27PcN35z9MCCSHJEMTzECHF4kIAhKC/alYEKshW
nWX0SUeUzBvtmoEFb4NSN2JQY5f5OnLjzcjQhVFF38mdQNutDPaqhmSa8LOnV7MV
teOeoRaeU5AC+0j4y6heJcPxnFLKRha9oaR1ZQkji+pDYJBwTBNREPt6hjY6IegS
L6Dxip3v3J9dSD5gOH+y9gInZcLhq6EpFQRqraEA+lAxJdM4oyHiI5EJreS0s/o/
FAt3Dy6hdyJrtriJYhjh1M3V8ysAevj0GUh/mL+7QEysVE1+L4ixhZNXURazK8Qn
Kow1JN+maZcyEAC2V2hw2LG/F4r9n8Mozk1tD/WJncGmfYdtjb7Z3ktei/vCnKlF
HgXeLxmV29hT85AnJiANCgps6Khj+ST1AQSMnpu16BntSGE7BlLZ5VKphPr7nODR
B4rd8TyLnD3aPAfDDROuv+J9plOHeURb8DqFKpthx88tTVPZ+YL9WV8+tYArBxGL
6sKjTVnt57vLb2nQbEXY4yzvrj9HQlGGhIZl+w0zZPdBH1dWYbyPI9gpmXTpJWbC
ReoSRqzDL76UHSNwr1jGJ3ATCyu0aL7DphVFtX9Drw3Y7QnKHJsV7bxFBF3C0rA5
RYny2n4ogNh/AwK6KpaFsoH+3o2Kt2EDL5OfsVFTLIqwGtVUQeJxeZpzR/uZJEyA
sA7IMRinjCFZTZeG6WBMQKzoyOPKae912d2qcAX0vktpxEHr0+DPvXUydDgUgYLs
f2K8o9cLmfM1TSDlNAswj1RIufBjZsNwdoe4uu8mHP2PTocvMPvrhcr3h3ZA3EHU
mZbuNAvkdOAmLOEBPOJdi6HkLUWPm8hN9vJoAcBk6kOP+LoQvC+QRfxiHfbVCfOA
DBa1ksJj5/MUCRcH26BtcLgluZDwmxtxcCTzL+8McPej9/V4JNc6nKBD/fxm+JGP
5Iw8wD159yWV+c+qWvkKvW57LUs0W1ujbDyRObZne4SeRlwv286lE15Ep833Bvw3
gv6YPos4ziHtS2YLE0ICbdnTSSZATVtT9OPWOu5Wrcj1q+pfBQ1P+f4O3CxKmuUj
ebtBuwy3eDqIhH0u0etDlad8t9BIrFXQ+NQ+6gMOBKRjEAldTWBaO36rOvlVQQUO
sfPUPdywIudDgi5QdJxGN6xnNgSY5hb2v4GC/S8TovXVzZ2FGYFwmKLmZbzZHsRG
ZtkuQSXssKW6aqPoctGiQ2tlumJa//F6elOS2stXGfB5OMSRS0cSdgNaoAeWPNPF
0clWG9ETHvLCjR9CLj2/Rn/hu7j9aNqcNMHKP91fUDML8Bif1dAPfrhsTvZ04F1W
PuPsUh5QMzr/SLKTyIsa2ErZ1wylSw9EGwJ4Y9QGqporrKSXAIKtayFqdQYTR/yd
M5w4zglyc9YbQ3YYdqw24wCoYSRFMeGRaXQH2Q4KoJJWhISJ8BlQooWJImLF3zl+
vXE34pgObJk/wQh9e3f+G7V2N9znlL6eHqTwdBbJSfeHFhzfZwxY5KeHy23gTqct
rgAC3VtwJmzJ7lpkVF61s8MfHxshuqQu7DBKoLwItC8XCmro3kfqs3rCu9Y2Z/mG
9hCjKlU4JZ00B48GZJev1LZQ+x+N4tLnoi4ozwHr8en1MlkplBPK2IVKeNAdHLV0
dA958cbKl5esaCyfwHSOE6d2EI847nUGEzLUeGI5GFi1A2zhd7jrIL+WXvhgrhqK
XhAOZ2mN9CHOx3VqP6IGIemwq1BDyc2Hmuup9wwR0cHSX7TjM2AmAOM+q45M8Pko
WJyNFUEM838X71/5ioOy5YAFhLrTgFXbK7ogPxy38h5wHEoW3uugJl3MiB00yKXi
THt5KMz3pxu/kbhwBow2sSWJ/LfZjQOWJd3bFh1yypW06Y28StTKm/n6SqvA8bgh
xoW14rrlT6nvo8t73djIbZrLc2pq9qn5cz9zYHmbVQc8EaB9yl2pqkxjF1UJOIk5
KiQIvwH/HvJi96Gg8HAJwERSOioumlpkPKPxSfjnijjhqpmuojAq0FPf1NUxjveN
oMMcAWo8UbFchHPStV9ZgSn8rrnkdcQuAOEVcY236DySEzZ0ZJy9Wvc9DXb7dDcc
8tgMfUXflxr/peT/v9CAeIMpWS+FZQKrnoUOe8vEuvbAU81yST22D8f6d9v77eG+
CmKVxUvqR34SIWawhev+74z9dxzV3Uo8rbayO8h8GF4sV9qsI0AlRzC7lZXCichG
ziESsU8Y7ui4juD/5EkX2uDD/B58Z4yhR3XtLxbl22hbVRVfmAI+1pq8M0JtcVB4
Y+ZbBXbVE9uIP2WHnNGCvyE+r9+7epXLI/BIdFY5/iF5GnIhwGS+OVk8DKbBSfsf
QXylgKSX/kIUeztb67AxYbjYVuAc8k7FlbYvNuZLW/E/9CbSSvS2AtEcioS6ww3z
ugu3DEnHg9DQZqS30NBnFncJxPidQnx931pcHT0F2hI21S0yt7CLd4V3+6/UiQEF
e8r8FL/06nEg07eHg2CB+1PijDpkulamDJzf4aOYAdnDBmqD7GT3fIHNXm+YK3sn
vfq+yTPe4cTKMBi20a5ux+/Yc/pk3Fn7TliAlLEsgER+Y4iuAkdJ7q8FtUpVYM/c
m1DnG8FN4ZtxSYuA6bFPw/ZoGOlKt4Isq/qR7xAzX0PDFDA3OUBbNY0pOzqRXLVV
M/xC/l1kjSWUWjSYx8CgLb4dxLKOqOza7C87Z8DKqaUFQiTo8V4ZzMNSKn6G6AmN
OfGs5waMMWG+bkEwODakxlwsIjTQSBcp9HODjoqeC3CezMIMWvvCBpdkr6DXgh29
y55zVFrZ5obnq8ZBXJXPcPJ48X9CRLHfyikH7KE212smTRKmW1po7BWGuU8r2itw
nFniaVLpoh+kbGzyr7g/H0vgfNKppsKkMBzG4pZKNWEDKDC7iWMcyPD9s+MbPC2m
Rrmp54ul/yT8Fogu1ngoBLJ9H5R22GB3nel63YDJ5Z75ARGwsFAjjPXQBp0KTrb3
9mnaj23eNic06u11/JInIZj7ripETUG0FncG2eD055e70lV5NcDWxVhs5ze+aCpt
OeLyW3E3X70jTMZYF0PhrLhF878u7Lpdy7puEe+4OGBhUcONTdYshsT8jJTfZuMK
6ZUnqRnt9kGY53wSP+CFlAhA4Q3vdBEOlXTVXSuhircsnBOreF+E7tZ46m6Bd1x9
yqwdEYV7Rb8CMxMgOgog/B9LJLEm298hHi4KTSPra8QMA0Ig4ZxZ43r2GTinLKph
ikOaozkmBiIf2630t1sqKy/dZ6h8eAU5T1XPETowOoEX3wuJq0tXMyR/jCpnZJLu
1aUjuFKTCfPW36YVo8Odyh7hTzz4FXs/drFXsZhuLFCDRnWSMNXlqOIbJtZJ/vkt
Ivw6GZLtqEj93TWpIIT1onJX2VWAwbrFmjUhlGO+ImdA9fJd4oLqiIvkaqpD2+nP
nOXATaMMgs7ZWQckYb4mEKB0Y2EUZItRg4RR/RIZljxhyqXh16/pXifp+a3586Gp
Y/kQ3SmhRZUCMyDhr3ovkOFK6f3/PjiwwIxKYZhQzya2mlZj2pWX7nskZ7wD/dU2
1yPF7x7w2CR5dxmnwWGLxUi8NKE2evjLYuiWXRHWRoH6r7ymPJTjVydxnGRqer+Q
45bUeIaf9Q0GB158IFUDWUM3puSTniAGOOdx8VpXYP6wVWiFXvcTSoT/ukm/f2ts
HCWgQai4tGXl35uCGUDL10zB/ddFcVl6WHIlbqYoDEaZY3ZFqZT3DntxrzXmilZL
16Kyi1DOjpa2ygEpntwRXGGJghvPiKOzaaReKxQnKzvvlMx8lFYYSC9XeAmShX7C
CqGFI35MLNyXhAdmWK2FYeg2fIbPbzkxzM1tUgS66R6+VpkA/ITz5HkfCE/YdBP4
fozB7FsKe+hgZ7ftpMvcP7CFVwnAlk3eDaftR6XSCvnTjA8WSLPLqxCMhTI3b5wT
sghi6thPz50AiIWQS8eVLjkI4jP3y6Mr42Vp1gJJYXGK4f4+5JMzMFCzg2HS2z/X
Ret5J4jg0pW7yvrGYmd7kcOHzsngEVfuy4Rlb0uLol0035n/y6kbOaGXKY4lGTkC
FAIk6yYXgXIAMqhWNClIiTwfmsqwjhtI6JDXMUY3FJ4acgffZNN+OOLNibKI3OvB
5DZ4y33pl61Oo6//56aaC8OYGXW6KBJCjLs1ZJREkJpI4NcM8+7SKAzS6O9r87j3
3MDAZ/EntO9tTqZEITZH63uLeCpH61ufUoCqjl3i69zMd6VyUZMJmY4V9UtSoDit
lLy9rS4KrK0EBmmZ2SNsLBdQauk85CM8790/n0q6bCVtje3wBvaMJTQQpOXdMtn8
qM09ywVBYHcd4AJ4hZYz3yyAwQJMVWmBtGSmVLtCeltpv6kYH9/9L84cSLlzVbqw
NynUcVvX/uBiiB8Z8fpYtSZQesLt+mBCCtDrPDh/GmT33KSCka5VLSj/bRDAR1KK
sQ2XMDomiGP4lbhiEXBuQt9c8LyEtL+Z5QsJ9AaFuKxvp8m2RKs8jadoBIjwOuel
i2G3EsvXTOL70cSnh36O33rdFcoUNB0fdgLgjCHHeYyPqGkc5reWd37fHqYRKVS2
vOO0wGHOYNuRkcnZOF/+Ur2H0IlM26CIOKcDXcplYFAbuX73PUA8afI8VFsHJZ3R
5+UO+ucSwGt9WmAe92KmWT+EdHbAG4apb5qvBUvqj26PiRFr2S0dVjFEz37c9wWx
tIdVuyLF6GS4RXK6AZPjz+Rsl5zEeanymxzvU8Lx6o6OrrJsXc/a6/A25VffU2Ja
TTTNN/GblZji0ng/ExToxdW72p/aPHiYUJ+a4NVaa/u0j6guAOStjZW3RPGz0Hl5
FOXdDKB2UXswPGecT63duXeeRE/46fgWIHkmol6wbsFu4f/L3jobCycgc1i6Ky2o
dgGmjELW7RiQPns339X2qytULqR3coFXVNJ6mRrtrUE1MHkpK4PuXRSZUTpzEZBf
U5sTyKWzhlwD1gGAF/6Mn19kv8opMqLvU95mwm4MBKUTYexcWD/USumaqTa6tUBk
boXRRpb7sHiA3RmLuRMaHOX/CWkhPCapI3Ovl+d8PDhWRes9GbTHOvS9Wa6fnbBM
t9vRGuaXetEzveGExAOzwlRByBUqHa5kvvm4udl9BCHvAPcJjc7U7vvVc1K84ltA
qbD9yCLZ/vaya0O1mHH6biaXrd3mBrm0qFg8lNtM0I9bgvCth05h968ajQSu4qY4
guuTDvx0o4lyzG2E/eFXqUZCEigVhf9+L5exaHgwMw0Ta3bTAvYeiQ0RGmePssmk
ShldQtV2lsp7ctlo5qUgAzlmo4naM5yqXBMNy79T0N3wlPhvjbX8610s9zDgAkpD
uZ+dkjq13xMtnIumVsAkG4UhxcwAMQ0MnJgncXuz2tt22MyHPkfE1MGwLLJqbylt
7X3ojCsmM9W97HpfODtGUowpHFh9uIhv0Sq+CXCdR2hnAJIt38tglr9CTT8zqqNt
d5AiKVOht5r41MT6f2lR7a6btiAkY/GxNNNvzDddoJfOFoyMpscR2IRKwZS3pBsN
HiZ14qGX2nhCaLRt8bw/BIhO+fWUl+kI7wLQ8oet2GbWZzfs5tUXV7qvTQQJbtV+
f+arZRtXPqvoA7MwpMvFKMFEPlY9CYNY2x8f1UgKdN05EKcZPSLRYVN1CoHNa53a
3huvcaugewqO733Kust5oSm29Zn1xuAVwweRBpcmJ2A4RsdcJUQb/lEyMDfOynnN
vORpsHcB3MtgrTGqGqX2l+uBi8yZyNy7ZsqobzJ80pT5vwyRiO5l2oMCDAFnJCeC
vUSkQiAc2cDSRS45PFj3Sb8k8j9Ijg6AraFQk+0wstok1uO3SwmEG3JSAWKgrl8T
5z/DmEc+TukKB9FVddzOY/miTM+BN1huwhRB0J9gvp0Rv2iv07fsx21cVa9sFBOB
Xg1evua8ZDYMJGGMVzsV8IsBg7LuhORkDYbA9AKhCzqSkBFsr/JB7SCVq5EImMVh
P2+wQRwf/DmuoUp3w0nWkerd63CG+un9iPJkan9o41PXXprPjPQ2XLSj8fhVsRUN
Y4/7t8wVhtc58mtfd5Jo8leoFa4Q9EuYD+w6rpH0b6lPjVbYB9KYHB0QG/27MZ7X
mhJuKr1ak9247efGi9ONnVlZfKKSsWZQdu4h3C7lZDNqtU3Dlq704TX2ppSaCzSB
U3cKrVzH2QlRHe0jBWJBhDptmO5oz9L6QgLqNpRnX8tEJyEb2c6yDniCLovhxPj9
QxOoSIINM+MIRGyhBe/m6stCJ4i8zXWnE8h7KwgKCDRLtYVYRXGnG4tkijWlSFPv
OWTBLHLdSY/9BlZw5/JstG31qZyzPASlKb8zkZ1jZtuCT+Oj4nH+eemGkSvIfpAi
PqYHf/tMCClRaadEI6L66JsMJK/tJ39lYqoBOL0BNon8Y7cdmmsUEzELY/PtEz6A
dzq9Qq0UzEfywCy3UX5CAlJx6+TrS3vRpEccflaBSxNLIvFhxTh/xnoZSdzi1wNy
YnrwpGxd9yNZ7AGq8rU800a1lDaTLuHFxNvRuEQpys/2GlHPkiWq0bqiC4VGNHum
74Arhe26CsBZrRpFerm+DuxJAXeLwXJcE1Ctz/+PIQxwwjbbtxfleUaG2Ou1zkgd
oAxRDOCxfKjuTFEtNPxmyzGJeCBXMtagOiQ7MHDrxJz5toQqGIik3+OGR6G5aY+7
u98oae1IQ8Egi6Tr0QjXfF7i2rbu2ttKWTA8BrpTAfgAzPjayLw50LE1aEuH5wN+
HUA1LL9XNkmTEW9KD+rqZMgbBU/DfsyP00AHP1cyCSpl90mxl5I2+xadlDzropV5
oAMT0fjnhvj9AnqQnSFyHbninpqjertc1zR80UPfzC8g9HdpfIdnDqfIDKuvZNN+
Ig+kVOAkvRIn7oeo5MgobrwpuFNQnBaAgTDwpHRzUH6ibR/GaEwAkZCaXfpADCH5
TXpwc5SBBnAeDMwcfp8GtdVJAtFQl8fHgJDuNUWI3n2jB08EwwXRvhgI5vlOr+Kf
HlGobhxRjOGHw7bRtoM4365WOV1Xpk1hR39nN4MvJb678OVSBE4zn+m1VW3kvqHb
CRH6xDQ0RtvVWvcVbPx2jWwMsbMEE6UJJTlA0n5vmM4MzoynkZgsAwan2/2Ofgki
7k/KO2wHppt/+oAugQCdpFFdJyp/8l9hC2bSLTyJKXzdxEQIbpBPqDVMIaDbMrFc
M8Dn2LbIXywTmgbhFxpSvCj/sIz6vsr7vC7kiSBSMsu/h3g4AuTtWz2X+L3j+tDC
GgmHC/pDF+2uN/DuKXqpksBOIcQltrXU7eN9wtgeBH9gC3HQxc1oJZ+5TUQR4mne
E7Osk1eVApbfTpHhW3Eeo6NbDVfkdKGSx6iRxwzSa82Xu0xTm3IzRztMJokTtsbF
Q2V+Uh5BHO4CpQ0C4hE7jT+sd5tis2POYycOME704JY6daO8SB2kGuZ7UlrNM8qt
y0Ri0bqM91vrTIzRfbsT9ClViKdQVQAVSbqV1O10Ry9H+JAVyvZHQdlpGYVSeEvi
pSwNweaa2KwUXuY6s69LPwOjFxzejO0QMRG3uG6pfAGvr7o+iWPyKwoS3O6UqIZh
dkJ+CVt5hkQ3XRy0dS4MfImuetg/BvzkaTgH5XSqmf9uKE6KW8bNdgUoBwUTb/RW
diTVLtqP8R+ZHgZ0qeaxoZLc1DK/sPZhqiroqW4PFNgTAUSxmDdL5/dnEp6y2oSQ
splvwUG3vTsfXw/PyJd3cNrFcQ4O/pE+H/uRhwk+xcRlfJGTs5u8/I9A3Ae0vk6a
Yrbh9ZWs7v2nUpi8XEHyDuQyYrCA/z4f4Efs6AYYLs1wo4Ro8jvY50Zm2+bIS3OS
Ac3GgpfP5wOpI9c4qn3sfsHPl8M+OUZNrjvA1iRobsiynIL1n745TJREqi+/WDP5
QkHRYV4GIHgwl8a7JUJRobW2kmMpuzE5jVdhhTbQ1XJmmwMWdTlUZDFZVdpuP5O/
G/hvSkrP9GHN7suZKR21HYus2O3LyIgDoohDBto7o5KBT0HWVQwmcIxEebyV5yOI
frQA+goy/ReUpZwgCSC/eydCkQU9tOFzsKmsyL2nEU5AEMVDmQ3cmeIjJinypgxW
PoiIOJ0qX9e5V5ILa564pQuxatu/MciQ74kRdezjadg10VC1Dc5HyzDNnyQnTn5j
0eCrJhlCyQTeni8YFylp3f53PgDLfdyvOh0DgfGUEGCCDGF12TCE4/V3zkV7VowZ
rDPp3ztbBDu/eAfww1OrDJ4gQtZ7D7uwGQa3JrftLAzLs44iEuU2wVWqE4CtAvjj
zXpeHvaWA/cYFpcgPdbDn93kCw3gVPDCAGbkt3wHUyRtwOzVU1CAzTCsdoGnQGtb
HnBQVModDC101eLMgig1Sw4ahksd8TZ4z0i5vYWUzuzVN/sQlfPIJbYlVEMFD/WN
bnzlOCpl/FnqKrOKPs48wqpoKxy1595SEUL7KtDim66oL3LtHZ65r9+7N0Ujf2Kc
xk7r/3sWL0MRtOZEgRRoXG/5LrKMpqG+wniK8Dnu762TuQAGGS8Jx9Co0BscxoPT
0Ek0ip1jrrCL4i/iUqBJlON8dakD3PkHwWbjdMANq9fKU2lMqhklYB+svIbeC/+v
OhJX+ORYyheCNZcaHwNc038iYmcurDv2eVw/ya4XEEaLbg55JJ5FErZLbQ3kYU8b
vmi56a1KP0AwT5oi8d2goIGL3RtdK7E5+QbWdGSD0aA+ACxPgNd7ebk6Jq8VHN+l
fp9xYm6YNFLqSx3aqRBbqmHlPcAT+f01+MnO+AV5YYb3rnCHeyNctXvpEopN2VvR
svPnq9az3wpfrvLaX12Pi3ITvMvaw6EmiOCfUvEPB94SrRwY3mXyQl+A12IJHl4p
hYbGVA/TKDL52TVigAOMQkvMvT4HANJ/KqSPhoQJZ5gX6Ybt+JTmCIqOU9XhAju4
xP74vrjxdkyvRe/LxVdmgG04o+/zKMV9I2hP5GlxSzMwk6tUXvgob6fCVKpY/uKr
EEC26b7AlVG1xI7RedXD5RKBg3nf4TmhkEoZip+FsGIb4ryeyP2HJv6YjxLdbpNV
6ZrpKXH56GYlxwPs3cpGFhYTAClrLLeB2mvdin3F8/6RxvQjjBvzlsfKZoyzL+L/
hxjgqnl2c4hEu0M2Ab1x9ZNhCm5bBsadAa6gwdrjjHXhwgqD8wEu51SirJw2XnbM
O4gXzM/oCWanUMqJzqoSAojwbLhXuafzaTZlnc0PfnR418AU6302e1KrsS7U+ySj
D6ItFfJdRa5YOqluxqwy6GD34PZ1RBWOJWexB2hochtclreflRCjZf2HDPHEvQzk
NrSksYl55NeeiDutSvKFThUKsKTHYVWAlWVswancRp5tSoS23hR6LbM4fme46yO7
D2O0OEmJXymiJTp3XQDSLER+SX8at6rQWqGsM+hfdhOR5RrR/zWSi58t7tZNRDtQ
u30EaiPVIGdYO6jStUN5oIqxGr6fZ+1DJ2Gu1kHhtlQa3X9n+UrB6dALWtarNvYj
Cxc67MOiVVXht6e6NvZ/8vYJA3PHj8GNEBxtd0mFvuANl/uFi5DjApmDoAImwjVD
coiIMJj0Y7KFqcEhRaWnPUGBeiDDyhxEFnG0Cswf9zKEKWN0blWl5QSQOLLH7dGW
LyUFfsvAn9oFqJqlzznm8TFKuTaPGi7kB3lLiadk3AGTYmGXFlQ1yR8Mp5ZkkxwO
wSRbQFaR/99BmtWIQoGXQ1cQg96Mg4aU/Z8sBFxoNK8IgRLJqYyxDsetmIlwzUsN
OALfpqx7LenlIUy04P2qR4XKFbSB2XZxPsdr28y27fVwGYzA811WbFovgIaBha4h
gi/oh+ygAF4HqjwkI8fmN265+ZqyVQix8ZRy9i7kl+66uYZdSlsqiS0JUMMs94iG
omwBuRYmCNVfquRKE/9C+Vri2AUxcC9V/x99qOxg6td64r19uJs/pdnQkAXwydBm
LQPfXsHU7RBQycG/n8Kg8/vBRRmFms+UcGEPK3hLwrypfezPNXUANF9Y+t/LQ4dO
doKGI2Vyh8Iu6V6aurqYPYjpbXkxrPGyULKk5mNxpZ7uI7ZSebtbkCJsS5oJaaWh
P8mSL5CyD3A/vPy7EbAzj2sRgKVypiAEe0B87WlsLfvmEoP8EFOJIzXoWiPUnYZB
P6VI3t81+tv78qk1K+hFy5QGO2/LYbSWpzchJOmb9vPWavu+8STRcQcu8mWsvfEc
NdZbnJi0+Lk+tDJ20UpjluR1LixNRP5wqUQukYUza+FbI/bkM2L5eHGcQ3WvW1jz
cWbxMrxtiY5YgnDjIWrjME/KhjqP3sMpXBLsp+8tKmt81gQ2MHTUDLIGphr9ePaL
FaDo21m0sdK/MB4w0zjXk8Ob2LngJxn2nD45LOaLenkXw2JgyYCzADfeO/sJsqHh
8A0P9YUup1sMRSM9LeLqMEkY150PbkEIbclGVARCzFBa8e37e66kRDaMG/S/Av/W
aJqy28J3Hb20ANMqYPBnjeLulQNpjqpCw7QS6hAKcPRWHf3vYB9nemqBgd1dmrUh
IQmyDMr78Z9R+S53vqQh0Iz5fCITtw6iaCWKn6ddPnCiZOreKt7ou7e0XXIrTwRS
YfaaXWw6fE7Q4hBtW0+rxS5PISJxGYNpN6RU/6boT0cs9g+UGc1UsuJBlrdk5hJn
w386mNCC83s/YavYKkqHR/3HzJz+NKhMzcQDhTxShLwp/lCThUEjw2pPfrX32ep8
3GqA3dtlvj41KK03IrTWphyvUT6480ZzUCrw5tu4wpNwRZXcYRZThyFzDwR7+y5+
XFG7QjajlCvO4vbLw3M5OD1VlnzbJbXiFc0CqlJvZks+tSDB8NL6mx8MY/hRQuGv
I92kjo48ow9LDYTg4ob3YzZNOrbrm4B7jdsiBRy9pytMjGLmrhYsIA0lk6pb6X9C
wcM45uOTqJgZVEhYl9S7m97rkjyVUqyPcjP1eNk2djHD1/X6Lk7PWvgW8OfwrAgn
dLt9PgnnM6Kqv942d8llnPLUhFkuRC+i4OOG/2sSLAFlpOKS1bsktjt5fX79ylpJ
lj5gxqlKNariMZVt1JpF/GS4ktoICGUFE/qMbb1lVXy70vRPRHSQCd1sEAvVnrdq
3QcMg6IUDpXe5lU8BS3Fa82pXD+ILhVSS3LME4tw7QrltV2bzCqKu5h1w8xP5sJ5
89z6eue8UXeQAHZgEVVHnNXH+y3kL3nao9dazjk3FrmdrXcUv1ReiMB0rDbekkF7
6iB80HrfBOOGPCsO7MggixwP8i60QuKA4byne1OXNkglKw2OR5xFErc1ijpZUvcI
+4OhVIO+qLnVtk7mfGI+NVLgMRenwDhzZAvYuXNt/3Xa++SSvbTVK9ezEtshEeHq
j1qQ2y9D0JIRakH10fj6B/mXK6RN4CrfTXcxpqs7GmBRq28rD7qbMLKaO7j3MCyN
ZnfdsKibS6oA88Y9aoCN31HXmdsx18toA2aySsQn9lq+mBtEJXKWNRW10/u3B4Os
Nhk0xSlWAQ4RUjWlbbppMLu5GYkqtkDqWzaA4fXDtY+KYVy4bd0Wp8L88erjYhoM
I4ZZvaV0BkaWL+ijpMjnfNd6aj4vREb4AAxxOlftbLZLlL64xwjQD/kkK6OCU4ms
jV2NJSFzO1ZW6ttpLSC7F1+DntH5uhOwIZwsMCVbqV2L8y/BeG7PQFH2oc0Flyac
aP97q107EMmN90K3tkdmZEA/yB+nico+ExQMHHDlFlDdW1u37xsprlmmZLmX5hN+
/eqqoezm2EdsEg3kinPsxMr9Oz9zxyy5ZKE279l/yilmVJcSTNQsfH4VBoO4VRE9
tFKgdwgfNA3kESDPzp8etvpclQnHwo68f96QcPSEEA4QRf/cNTfLlgW2+ZPU50a/
kQjgEzOaCSKKzn05mx4r4wyKTk73UExfHt6ECiBX58djCsc3lyC1m+Ps6AsRNuaX
fkuu2y8iuRHLoN6OeeBL0URAWf8cOLrGCo+Qk8vIPIPYti2mTcjomYkCZnDIDspk
X/ToYXxHDeXhyY/yQWicaYhbolZVUanfRR+30OEB3bP+awrqEH0KQoVjYKuc6q51
fiNmYqSijIyDA2s6Yf8xJtKF/6N2t7dYEk0p0iURa4pdCmaNg3rsymk2Yd+cU69q
mKFtAhROWLdR6TT/5CVwzTazQbNjdz1jrqeIWeGMIOQsyhhRBOzB2WmVz/G3W+gi
tGH03ANcu+Qc32jZpPoNoAi/VtSjnbO70049PfU71nI6+xtW2rwTNGQotzaBrVTw
YnlGIbvByluUobBOZg5upDMw+Vz5LVht3p6Zm+Ob8xbrAsvP0ftdr/tMlQXm5eVv
Js7X+ZIExr64ahnyOSQVV9I3k4WPpNXQTnVchcJM/3fexF2i53sQGINAEvNaerCc
u7yR2ph/UDo44GBxZa8FX+1uaT5oFZovzVK3EBOdgMirzq15wAD5lMZwnimpPos0
+Kk4Uz0rgY04QSK6i/72v1JsQRB+M8De1U0St9BhmqJ3RwsIaSXBld6EMuYG/SKE
mrpaDsXSdIBbs9Hp8czZjAxABythQee3hnLj9kLwRAB3BsBYr1zau/4KUY3xJzUZ
et7DrhGDAartD3mKniidyyLdetUiw2mQw15q9A2KGglGyVEnOJnWxBPX/lVd3tH1
gCPgGvAyHL1CeP6HaXV+fMs5gFBNPmDRIH2SQOk44up+Nr4IqVzb0QvfLE0tQTEX
urwfUqrTrDT4qEgw/S15l5lXW+Fk9DsIBqhyWylnxgMjKAge7zLLbSObQd+Dw/8u
d/sp1woVMVnUNT6kwTOBq6yMQIcr3FnDBhU7n2BDIEZ5uUKQk0O/LDSexnAXW1V0
bWQ5C7glaRMMTkdrNvYHWHgI6qiBWjis2kGVCch1/1ZsHAtlQrwGf7tlDlxwzhIR
uUzlYp+Fyt9/EqtEfBW/lgOb9foAmT+iYR3TW8/iFdHBBTmBkcCnLYVfcSD+BgjT
46MxGY0c1DfNuR8LFFvIYAaPdCA2CC6DeMb3enOzD/32NYU+r2MGD5Foe1qp7+J4
mFzjplg5NImejSioudCK/YYZeF1HkKriixZzZkKjNPd6BpoxtuGpaM3F65uAV5Xr
F91uGRc8PqxNEw+SskTUuixVP3LejZ1vU/OHdbro/4uAMJLSFS+W2H9IN4V4pHi/
o+VpAqpuHVXIxKREo9KkiDz6XgaE8y1mUA734W9iVvvRsgWfcJxUXZERpjQT6vGN
54d46y7E42lXDYMumeivOhdbngostWzY2OSH+DYO387tIYIlK5uqbhaydgsnmLAO
4dg7E3610ZVhlW9Tcwg8ZLgpdYnPnBmx1JUZ0TvIRywU+Ja2WdFP1tMPT6L/vkFw
Eq/WGuw4A9mX7mee1b2G8oytlPWNcB7SgIXRRd+aG6zaaoDB2bd5fKxNqKPNdafS
zC5+3ELhrWsjmy5e3qOViFZy5ZEgOSG/E8Sj0+aVJSLD67Moki28nKaddUijGr8M
t0vB8pV3gtx0Ysb7QSLLz16TeWrwopdKMagCNQJj427f2dXV/eymjUbArEgl9BiG
/vjM8zf7JugDO6sB8X9ltpyAEWk+PAE1FcwARcceqk28UKeGdLZ/V5bGNvsKHvAq
MvOpea6sQCkv0QOU2NBLeUf0F+w6nJwOLylsNVWWRFaAPdQzlDhNmr1aI+jz7UFg
4cSjE87pb6NE37gTMcek0RCADBw69EbdELWcqB3o/xBP+V2uP2Cg6cElGTrxoei3
PMRYRjIapI3K4fbnljEar+nC5bMNK6QPl4q4DMVqLFL3cM6l2ywKJ7KLLMYte3Qv
LAGRlc+4CUpWq8cS/CBZ8yIFSFvPZmd23NEKEBc0lIkfJdQpSZrrfE243g6gh/mG
o/XfQ8WO0R8x673jEfWpiq2g9YUXL/zqa/K6GJXtbemDAB9Sp/xIFxAWCnrZr2f0
Idf2/OHCFoHuj9fZW8UBINmcYi1oNrX/yUNf5eqVoM6Y2lc34W74gtputBcOOo9B
YjvebDIB+HTBsKDOSX9D9zgzW7XXFRillpxmQEwh9sJxnw5xTBVgc7G/KIMsKmbS
Xj9zDNFS3kIVv5i+Yl4hCB49/xqTRtNBVFmlWcaWPoTj6Ql5lbYVfG0LkgLVxmMa
AbwkKHUWP8vxnxJCj83SKC+S9BkjI9j/isWJlN6FHc3cVbA6oPZ5rWaUmh3GbuMD
BEiwFam0NOJMgccht65Ku/OiRlHpfuhiLfpnVrEZpEK/6X2jvELb8W5i22NyHXYy
nO0Bt3IVi1GpNiTIv4iRjF2z3s2/ahwbnkGC9YcX29h/V1S5NfKXzApKiBn5JafX
KaA30apeA83oAc+43RzbEzfXKyPMK60fS7D1LTv9FVu0iJS7qpkrlgEJ4zPM9RUP
Ms74MexY3JdBzuOLSnZ1K0eXmURfTdOk+U2ufj9h8FucLiKh6mj4lKnCwOMkzsEN
iOns5J6Q8A5mAXGInKCYCwxI3YcBsTW0WDvvym4WniENpl2V75tFjTRnomYnf8yU
7VBl+BRaVEooTXFa6QACQx7n4tCm+U3ZQGTNmVa+UbCukUVp4/B+1Qis66I6AwC/
ZtFAoklgTALozRT+DnFHYMercBCC3qjarTr1RIq+lpJnLGwbF5P4DLpdxg+7IqPl
WJqJoS8DRy135REU1u5TR4l4+AD+vdkcCX7cKSn6pqxJv8TBlJMGo8byq3S6XGCA
SJ+aacJCSe0DB9fdYE6lZtjh3+3HIN3A/fsYkZr1NmX5++G47KBG5CMB/IfuTD70
oJIFRTTJWBGMh/lPut4f+6B4CuITN3iuTLnauWEGJk8cNsREFJ+rRJNTKjeQNSnE
T6e90iWxp75c0hiegY7+OSqBCepe0q1apx8oxTuGzWBqBPdJ1nHw5b6RZkNHLuK4
+pxL4A9e4HD4/3/MM5+RFeIFbAKO9d5DcfhFnBftzLiFewfF8TXySISrogI+fc1D
CScn2X0wr9luIqMOkhH0msMY69fMSWbs9QBXwZO2mRRa3f4F7oZNJHjDmfsBq7RH
+49vYYF4O+0sm62Zd+A8VyDua51k2mlB++P/vhNcKFzWWexvs8jWa2+j6vsPxAxW
2EtT8/nlYCoMwcyy2vJiG8k7qEiQQN/UrTUz+pPsOP5vvsXJNlkOU2MI5FJ0AETW
vQ4TAGYbe1q4vJg0LDuxQmYWchjsMboxujebKaWxBUECUJj5cjSPsnRCK4zboXlS
PqJ1/0hX7ueaLLjzrYeK0ez4IMA+Sl0k0/d64SIA/Shjx7eWJ/aG3KtX4VGjk2IS
nZ+PHlI22pCxVTof59wGhwqeLbheWSYRMRcIBtO/DMQiAWIlBwOucHFjaY6pE4sB
icKqSrRJTL0DCnLoZcd+J+N23EsDk4SXXgllZKHCwr2+cEh0ULsW8Nxz3Cyy8cO+
/G4SxwXS2oulDeg4nEY2QOQqQbpbtBqLDN3WiBMLsEu2wOpX76FU24VEIOH7eNiu
ROgcjQQ0z1EsWAX/8lLxKeGq12Skf4zwLRvMWZm4sxY6iThneex4pHRKvVCS8rqD
ufLyAoJ8hOlTOpjuF0OqYWeemwsEmzZKFCDN2xySD4sfRB2rtQHCd14wq+ffS33B
qCKUIKG5UC/lGCi4cE2GQdqz7/lSrmL1ufzKuzhkfbKMbHxBbS9MzrJk4o6uJaYD
HHekAagY4KSQj6YQCHG1EG1BlTk3z/WXvD+BhGbRZP/dvUVfN5j1wyszEtQo1JpD
ovdCCoyNmyBmVdiGNzcAQ+e7z+ANASWmloMQrTI8VelAykMFOr4m0gcNvDeXLOln
BfFKSbeV1UQ7xSFZ4ao1PBd+c7tr5WXb23Kl1SJOEOtshx5OoxRNq/GoQHvgKY0T
nD07WOOSRTHpptXxVBkfsEx8EqUbo1rX0NhJ+49bUgDezZGmYmMgcAPl1CMUwiOG
vEPIofRnuoQQiVOLO42rNctpS3yduE7OCQpjGsTwnCShIUSJomcmOztzYxcDnkOT
2tVrJ0rl2CMNXH4bUD3QtvsylbBx6/3ct9ttNKyb2dZ4PyuTYfJm0QGgh/+I1Ea2
EfDEVVACy8fSHlVs8sSf7Dpf8USawqpwbQoVBlDCBG7Vl6eGUqt3HbxZgAkMBoqn
2o1iyuMawMNaI4RoupmdspnW6lqdUWOSWaVKXW0QRo1sqJ3SzbuGRp2H9BlyNBTY
C6xrgKyGt9Tg+osQtqwnuPNK0MeD8xvPpIjVXzH8hWjbbYap9dOWfs7pdQzxl0KI
p6YEAfoon8P2D+NKAHhfj7zIRt9EB/hqFWfs5qBgIsr6ddq7nsxK1AJRztT+3N4x
eRFFTWzW5ChF6UL/Soigcqn9ywkbEpYxveEo2jT5X30SKjKsMzSOxcl7cpWDlW4G
/Op2FYPRVeV2DBa6ftTgJ4/KNw7iMuqa2GceZXf94toqRHPFNTOsqj3j3s7mdIkf
3E9hky9ohN93fXPmjlYuAWNh700kDfVNNme2YT4YpnVlbRKqZ6Pdxs3D+L4hJk8a
aleGtUvHg12ecCq4OcoQsCXN/+2+cJ7ALTT61VWQC7TSjGr4uyvkAL6DF4uR2eQt
/E6XXWE3AIoNwGW7tOV7LpsgiSCSWoiKcKd3iUDq+JvMwf8fRqjdohuvxs3wJKdX
mMLYAAJAzb+yXDBDNHm8q9/QCSdOM3sT9+K7g0ki2s+BHnp0woRs2Krf3L4BewiW
SuLz9saN/t9NmfzGqvHxSM/lDytuLfW2PHujNhu69IbPM2GQ2pDBJndSQw9ENppr
SbvK8sPpZYD7XXumtcnyIm9J/KEjNUyvZ6fQ0KTWJ7qDcyAu2ajqiGhzM6SpD7ex
/962nYN2l8Aweir8Zo82TX1Yed05hAJy/PrDcFrRFyQF67t2bOOvUaZzCJkKolK0
GJrNuNF1BMHwLsCM6sPOPs9FPHDvvwVpexEBPWX/wIl9tLgYqAA3w8KESCi+C6cM
MiUDLWaVWkSrYGt4dNS4cctIUmk6gDJ7dTWKp46Np34yPtxdvk8d6qCY7tfKM0Sz
9lr4xpNBkw4vP5p2abQhOknpA08sE3Lx9zVwy4yU3jfgbVLyXeR/ryAfpvWi9QGN
vHbGvETFi2pB02a3qMyXzELjlR7YpjBzES+W0SxSQa6TDQl1n1fd3RkOQyGV0bYu
AoglRx6PNRf8qBCUgl8XHTJQ7yyLP8SV02IZ6b9phSRpEKgfsf3AiiEskDj6iDSs
/OIvdGDqcqEVgOL3BRnVYQnOe/SMdbnszfk977UQsXuMrNAi/iwETJMDY6tgbD/t
0kGrThlTcxO1K0cbUoqAQIoxcNsdd3GmBBdbQd4X0IpmGBrYVRZROv5S7M9DYr7I
jGDzBUZVZpxY2I3lPqgaItK7TC2w/2Lqtt0/wo7OlSwXz/QOad9tdmMM0cTaih7f
YO7nA99uPTxY/7XENSR6GYXUUobbdJcFzUvSVLfo3afXKpeWIY2vn9y1WZ9XxIW5
93NCjf06cNwt0q9QeHBPcofVaPjaN5CeYhht2tfztH8re6Ic6Pxk4vpCkVxBkriW
IZLWGQyfgsqd82C0u+oO0Banrk5QjQC8wfyJ7vnTn13a3E/rD5C5bR4B81/VOV3n
0iJOGUVJbxXl3V+feFZ3PRcKvyPgWcV17Z1CmwTdcanxz33ccfx5opuR0mxFfLG+
ScTEUmI/JUEhRg5lWKXbG6MjEyUGWpuxnZO+bxD4x9iQzkOciWb7oOvjurvAWGnT
H7AbrjK8vefmOpdD94EQdzobAdFxKf/JY44UxCjX5UQ56J1wq0UL0oEIVPgsUgjt
Hgozi8BhdTC3DgL2E94JlMN8O9ilWQc75ar14hN2xnL4Vw2AzuMhjxwFliE71mav
aiZ5hy/q3ixq8ggRaQoQVa99Dy1RDCbyvske9/CLHzgP7BIUK7yScTD7riSmpVoN
A6hWW04XVzMbETZPcAfkToquRPsPViiocIuSJ8Ur24ydre+t3uq1GHe+54JvgyCe
jMhPihbxpRdj57fLRde6KUUXF1QfDZcQTFcdml1XUUHruM9eMpMeNt7GpnGNfzpT
cQW+3H+/96knfluskJEWs/v/fw8g2WTJvLAvCRvvEqWrBkSY2+NH+nXQnwkhP3zJ
wuVWRuT0paPh5tFjOzeEISSmXi+xshyL2BainnorZlcsPGirjKy1wsp7ujawLySx
15NxxzA06pc1ES4NQcDG8Y/fBcXTujK0AE3ZPcSmDEKkwwxTkToxllrVtV5XsetS
huqnikdCjPVXflAKbSMvet9N8n8Kfw1TisSCKlxusLNceO/cIRpTfRodgyxB4HZU
+Q2Xiyz0hQngSz4s69h2flWkMYUYyGrdlSxiWLzgWNxo43jmTUhpAcURpzLs2uuF
re/UQuz91D/9efBOyGEPoC9Dq7qTD2zJ3WLdqhIiYYx8pQAbI60R6ht5zcjnBluj
5uM3T1ZzXgJ5XBb1Nn+8Ili4H2DqT9llvCAyEOG07lQJgd0+ub4RClnoznwa2iJe
9MGmK/qr2OuEqg+miRwg1PKp3GAYO8eiQAbR/gtdLRpDm89QDeilbr2CliQkoI+2
R2wR8XyeRJ7B6mv7m/DP4xC2bYzFLPYKU3iEilzFw39NVxUz9Hdsb5am6l96vMtZ
ARb/+P+aJ/NZWit/p9Th43XThq+WjzIse+8+803VJLMj48NnQIIOoqVBXwUVywd8
ewIG8szrD6ldfz1qEOabThJpavn8Hx9u7up4XZzBA/ukZSlc7Qs/AEzyUGVPCxZR
J1+pNdkVJq1W5htqRUhMlOWoZbpq3agmxmqaYCPUZje5OiK83aqK8Neuhhg/RlN4
L+NCtEhlKEEXp2nNaPgKhYTuJZwrlRF1yTlQkS9W8ITyXVIcLv//B0ju9fUQ5GLJ
hfdYaJRXEOhNW+5se5IiuY2QCvm3lg3GCrNcWqvsAh2pdWB/5zRCkJRpKCYZE6ff
Um3C9Bf+zHUFt7gKUPpPACFV8Pa3lp6ZUmnz4QS17fCNaJAAz0dk1kRsjWRpih8l
RbxeNc31IGKvAavtysPXPyGzxYjrZ0nrunIMIq6rcvXpxrebk6cb17roG2F+Q2/H
jmuA+jX1JjufzlwZxwOADXU0XsQDPuwX/EfY7iwUd6+RLEnejDUk0LfO9SqEGFEQ
Bd3K//f1nAdoc3KDt6YqpRPzUDAixd/olQEQNuti1YGNQdRzpICM9eTTPjNkbT4i
OjUXHGroFMlDJwyClHWhQYIoe3Ayg7b/DZJq+i1HH1ikranvv20vjHyUmzhZsN/t
UJy+T4rF6dqbTqCtTpK+5pPzFAiDsHt60+Y2Ye17nzEmH3Mjzfk8BcbAcZvz0Pwi
e2KUo+uOBdS2EQQhfO7iNZ/mkxJOQJ6H0bih2NqDn3JIN9Wyft7BmYTJSltMdWzw
cWdkLJvpGyctjxS9FFLqTlJO5OQbOcv8IdYiIDu6IL2d1/TaxnowAAGadaS+EYCC
ZDE4YGCFEKw71A3E9cgoeWSPpLZvvsNTBbUsOLgJ7ne+AHk45x3z+9SEdFgJPKEE
7tapvaS2/hD7NWXZnUVDUCrqYwSh8nkDCXACvlqnQ3s4vlxHR4Dikefio8j1DZ1I
ZQgqBxrVoTg4jNlK+KS9+OAU8xPD90ZElabuSCEGfs4Vw+wgu4cBGrgKbCc05OOB
naiLh+IAsGOoQNqRWPI+iOVuNzDkdy5ibpBEErXLfc00DvNfQXpzWYjZ3E7kxiuF
xM3zee8QC7ZaaiWRDZJC5RtsPy8MdDrlP4+/Dd24R9jcCEkniDkouiPx6B1UNwaq
w01453lor6m7o8KkPXtT49QpcpzuEihRRCGPTStSV46eWNVGYt5w+y1OO2d9RKgS
JbzZc+Qwa1BC/6D+jAmChg9jIfm20bdak1LGQKXDC6/NDukk9X4HUiP7xzUbGFxl
Y/sJ8UwNB9IXJjU+rv3oXAbUQhJM27KQxfAHWn/jULwTbh33JbvJTCyG5BH1TAjl
tVnyg+fsL5EIdH3odJnzKV5eKc1OVf6F18qrcyA1xW778VhaTljez5FB/wKv9WcN
tOxISofNYPsdaTKvY+56CJNdWPOF+XLNjTas6R+kRCobsqR/dO22PeZgMwpN5Atr
mhJone7KSXcjGRP567zFWWRMWmgsiM7J3XUmONgdC3hZ8VMRq0/G4386TbXXi227
RcOFD2ldASGH4fDg1yuGA2bqYy3pXHFwEf2YEAM7Dw3LAohA7344uM72xV9k2u9U
QP33IbygintKm/eHG4wCirIqivNE2otVamI8Vn4Vvft3/aKt2A9VDgxdL83hTK2P
25WR+DGYpLwqD1C3KwR2SYsa0ZxI65mFLApZmMeo2GuRq+Rq92qcuk5r+18sSVlu
KCcOeuLjXmyz0tHFSnFtgzJliOTMYz4l845NW2QKehwkEoPQSCNxWjOFx3DQOiVi
ljt5+vdefaAlO0dwPwmBqRXDfoBzDIHmaIfzBAAIdEZUGtar0F7lYcJKqunvEd8t
Q6vvAPohfwfeFB6RFgxHw5K+5L0QRbGNeXgCsGy5rDPk68eLYTk1gZTHq83LmsTe
0m+IEn3kwI6GSmW3BUTdH1TJiF79FHfd+Po3EDhNY7UPvMYZ65uIj7NEmiFx+Huz
a+mVNXZYFXeeMNdG6s16wuzDkDa+fuKEyvi8KrukBBYa+qCoWtMuyS7imLFT4CaX
LHOW1vhXe8m1BnSFMpPhx1B6lb2WJpnfnPnPE3DpLH4akB8wXWuvG/JpQ65Sex8l
9bTmQdnT0FKw32ONfqXu0VMK3P8Z0g7En+zGHRObTZylRzZasil05sT/Lta71SVk
mmMWV3TwPbRF1ofwcPyzuP0i3OaMMzFHoFG8Dw6whCwKLX3LHpaDO4WbFFjFWf4B
9Mrv9+n17ycqmdaWdvzTKEMcMZbVvRVrz1zHFqeTAZqxrZGnZY5eod0obVCCQtUE
729wccxtORwCxJXkGutgk+WMkyYesjXyjrc5Y0nswEDB/cFBLP7nQempBZPxoUQW
3yY25JX25M1kdhLuHjsInRUvvOMqrObCejvG4dkHUqdmdOjx2QRHBQmllceh1Up1
tkH0qIuLzsiTJ+GIjwNBI/LWl7troGcKhkhUZ3nzpCuYgRKrlHPjPjQ/SV3qFtHg
g5476hCpkYgQytC4392u/+4JdNVfFDLeTlJxgPUrIUKLdZplMzHcHqqA6/+Uy0jg
OluqgsWsyjesk0DxVl67PmVdt5VAjOvUmiRLMUxu9OKulkOyE7ObhpfD0xeDXkaT
Sn2Q/CiQLGe6HuZ9Xp18BMQWkNRUjW1GgLq4a/0esWA8YsLYPwdHbYQdNkv/g6/9
un50Jg2Ioru8TBWT3FFy2vkWGGiAJAJZu27ur7zBSoNwwSAQxtEjgn1tZ+WbVDNa
MQhkqTe505aA1SRotW+yF92YqH1GA0c3Fq6RrV/ntB7gLC/oD1ZgdehReejD7Z2e
J0xIvjsDeKMDDfqb7FdwDg90xm8bGvUZS8sl5l8N8/T9lDf+xEw54pfIbBCWIS3u
fpoITnipECTQzCjZvPv39FisCCuGAqkEwP3P1zw6yLled7GyZQerjvrWI+QcJEq6
6T0kQVllU2Mo8OtdVaRzSh/IJgVC1EnozgqX9Ms9CxZ6mTtbFwB4+qdYxFbMTzTh
fTfDiOmWUgdW6mxvU9EyIGsSpDpVgKYsQMxMRICrX1YQQoOp6vKJHTI6oIzQ50Q/
02hteFEuKAcCxXjIWW/fyFCD8cHb/uPCGdFsldDsDqSrWKq7owm7iRytE85OZr52
IxJyt3q515ZDE6L5qC7O+R21+t7FRAZw1O8W2ZbB9AaXv/p/uET20bkr+aS1Vtqo
g83Gcz/HUVFTeyFHBsnD5eLveUD+aeUkoFVfjYDPdDvK/Vuel7BmVVDutX5AhjZX
A3PMalJwEy+mKqg7n0vHdSrt35etYAvx+KIeKIU9UOAiD9zHZxOu3NfHTRxtVjB3
dZFTK5w17rraTgcXe7DvSwHbB9bi99sxUrD15hcqvvy1PrXH+RUDLzZ6kqLi+LKK
ZqUlnhVZiqdsvqjO/HWuDa8P9Do3fcIN+XSuD22eTGqiVq88d5DhI1q2FuEtIk7G
iQkM7vpW07wU+tHKdwPpJ92AdYGRUScyWt/hJDoCadsaK6OiXMgHQis+HtknwM3Y
GmGybXwFMbahEod7Alqwn3Ilf7Gt7jycA9a9dfqunFQjC7urjJen1GuDNp9F0B8T
xYn8812QT8T9OVhlBVQwPI3RY6zQbv/spa49md5YGLHO40gYuwhFuAFnk9mo+fKJ
XS9PftOG8E6rwvfRpoyH+pRT3iWLwX6nQ0iZC0kSRpunN0mNh6DJ//pnfKP2xBZM
xwvB5grYgvkU4pFiXy18l1+zNc9PYACz0gs3uW8AJA+jZAsYTP1E//DRMN46yd2R
HLvTSckn3yr0lHCmtif4LQCh6UTh+omw0MlsnD02cS6bh6qrUVVK2HDn9aWSe1y+
aiTs3oduB1gVtG1a90FabAmoWZjAh/JrMZpkd9MWDW6mm92md0KeU3JqX3cQZY8x
aOeFLmglQK/32KbRSjHxgi5miViVbYV0w7r2LkroXq4agIY0vupQRUqIpXMTiTWZ
XcNDH0IQwEghht+DHt4AMkyzmWXRQRXHyg9Rm1NT7mJsfKs9P0y1J+KxKG5chGem
HNgX4ucaJwib4mGfxiGuGetGwfuVkCGw0MwY4wvfcP4pZjPYTlAteca0T/rx2sFN
9qEUop+B/XpvKNJ3qTT1kleDnbQcDm57btvC37az3RUrKMRVb5yuMKf0AZKEt+QW
FQHE0bCnjD8kBz64oxkfSK/YE8xZZ9pkfQgGDhU7YbIf3HISew6x0tShGjHjFuDG
6crNMeCo7eik3grEyR6yxEmEJ6sq4ostKI5/znPjdcxWVVlHFSW6YlZAYbctDB4G
x4u+F869HdLzYtDFrqtrRe7wbuCbMVTtwMuZ6ecNgtLdU4Sp8hLbmw0VntnGEhXU
pmJStE/l6E/7otcftxoc5UFrwYwQBLbZ/sMNWL215VfQ2/W89FIdJ4ip7aPtzEfU
Fi0ggewACEfgh6QYCpaMgBO82K7/LRXdLq+9l5P0mmmpNUWqYCXa/AtuRHDHQnRl
67qS89bfU8NmOoQI6hUoNoimVFFFPdO4C7ag7plv7KIvjbntA8Jrg8Fta+j97vyA
uELQ23EH27PksBA65Yr1kaAyNpLlV+T2154ND8vXJiL+CczjaRarvwo0/1Kg89N8
3D7bDqhkbb5HIQBxUAvcEUVf9cdxGNwq9NgthrQWlsH0n9AP/JEMUMJH3v0X0yxK
iy9souyvTE/3AAc6kskdcfzzdaoVLf3tWV/lG5WO8bZ0nPWSqVhWADywiLzDVtCO
5KI+Yk118uqSnetOYqj0MKYgGN6jZPzU7K08L3sjAdhpeSTIzifujfxSLN9ApIQs
E/3qdtD+fNy9kIq1oXnQsFRve+qELGjTwkTNMi1EkfB/OkjLAj2yRC6NAaHu9KuW
+BfMR90RyvSQyrt1D/oytXA72sgMMwMZo5+Dox5n3ianY4M5Y0h5S4Dkms8jkVp0
GRn8ay+kWg0U6WQChni8onre1tso3CxBIcx2Tmilc5lmmECIaveFLql/hkR/xQvf
g0UNqUjESrhdQK22nKgnEvO2YoqAprVtpN7CstzCfDt5p8yGptKZLDq/w5tXijKp
HcRFfRkTEvfvQlPmETEUCzy69Lo0XUI2JRwrPAB/Fnz0F17rXGMMsi++1PoyDkCx
QO+NKvreMpT1O7josi2ZbyA7F4FQDosLZP9KfVx6lNZqFvaYAyFwALv7HkslGx7n
g3aw/ictocvS0g+0x8cxpOd5aMTCbNJcsKC2vli2UfjO2JF/NbSIzsAiJ3H3zZ9/
B6FtJrjh2OCCy/hfaR8ywvhpWIWwYe8fo6k4Ykf1EwpLDMNdzMWF2Vrf4wZexpoY
azNtupsSItDncFGA5VXtcGiwtkpXyP9kodKaUdYIiuf1W01Yqp9W8mV7Ee7WiBO9
GLcO32kwHqXMdg/SKz1DoxiuGpLKJK8tJHs6bsWNJIVv8RTDo5vUoAtNUn06frIV
jpuqSiCswFJNOZ4A6O8ep60d65W/PK2qvpJUuyOskicT4QCohl8+JUHItN5QMj0j
aemgOG7xER2xyrTMgGhzPfav1LN4zi03FH0PdUytHP/q8sxsh3olgu6kdqNSwihq
gus4vTN7tKvysmLWSdySKhTSK61gQQ5z4ZvtesNCR3KuqvDwdlBIuZtWKi+2QyeX
YHyyySHxakkJJEsv9G1YlKhRqhX/BGiKiJDs5Nrqf/hrlBy2rApIlm4Y9dM18o29
KqD9+joaYMwQFtHSM/WNJRN9Tnxy3+reu99rq4vSPz8mmChHMZlkNVM4gs21su4o
01GH4Sgg6/ZsiMds9GIZQgAaNnD05QUeRVDX7GT9d/uhKQPimU3qPvdOJKf90OF+
Wbjj4LrTmcLzXYlK6B5Hl8bTxstkO1eapxkw1gOtZCd2z0JGLiDCsTHMkaHJa07h
/lo8wLYTMSrB62/i0hoSgZw8JLhP/hXcSw0S1Ie03DLdNbdPJ8MX+09qe9vqiY/R
1n37eSe2uC4g7c8Hbl2TKmxB7f8yk2ldatDZjI/fyX34axhXu3ofxob8QVfOaueA
PDK0ZEl48JiCC3v/rCnFHRAzpunt3+y0uuZkGa08afqiySfnCAFDsEZg781h7fYI
UhzBXL0gt/a2VvbYknIt6GyFwBOyoKKZishK5zx0ZgInYfXDDVdXZOYhn372Bp8d
vmvy/8c02kMzdMIYEn8TDSgZjYELJ5120sFs4ZTVheiFCAX+aQcYOll/U6yQ7pv8
OnBtUCTR0HOh54h2MLN0pN/tlHUByzDVLtyjTjDmZnm0+PsM510TaOfVAawmzZjs
uE3aPUoYz9X7gtpSd11XNGmXKxi1Icd8oLQdag5+uCVZM2UBdNVdA396D8LMjChh
o5vI9GqWPWDCPtZcYlk2Xt2iW82TlbiGcvG2jOWRJhPHmnomDnYR8cbSCY5ftUqX
yM3dZTnVVNNna6rG2pLwI14cjaSTIBkKAYqZ9m/pWMLitSgNQ0ZSwmvnklfK6O7p
9jW3w0Ncd8G6kpeY8YYl7jzoPCZ5Yjvl/QwQ4ZxkKZbDK1QUkCuEHDdLKEhGkN/F
bNh2iHSMZBgdYQjGtHudZW4WL1qh7o9eirJHN/KlHOsmzFeFuAtOxHPoUtGk8z18
FJ9uv+2gJ/swRYX6ek30IQ9cszulXkWGs15IevGJFE4O67CMgQm3hI2geovzgpZR
nWQE39pjrP+V/veSyrPeFY87GHom9y3IFU8ljk1VBYk5d7gjmpQLNs32dEISixF8
CAhF6SRBlDg3qCk8fAZOXkKbozj8uLCsTkDosYC3iIJ3rY+nSTpAHc2uNb0eiI2+
rRlfU/5mqcF3bAAj2k9orlyJGJwAKUBrJY9fmg2XRlzSvDPmbpkcbm3qUP5FCfxB
MmdXoA2e1qClc6Yn1nob7kR/Qzb0LKjywym5Ac7DAt3wucZV7KtTO4n7SpuiW5kQ
ShZr31o54Ytb36kifJlNRry73PmiIXINoxXhMj7fnfrRc+LWWizKlo16vkA9Im3L
c4WKprEzN0bt6A4BEq/yGeC4LkQ25Bg3WRKNrmQsbMZoRX9BvsVN1LMDIcZWOQ45
WzlJwSbl5LzC42QbUzd3vWPSMtPnzEHzUEeYvaHv45nmMNrcjwwMCXDcsO5+XAAM
NE7RBCjd6QXWagxjwPsfTE0tJQitT+2IbTEKK1q4O4cEuDWw8M21L/tmf8P1v1xc
xGqaeFW/Lf9mh7x0B8MG1jA5natuVH15m4sox7o39S7xjifNwJ/1ONpH2oMmzc+m
tlGTH6RWs4eq5ViU/Te2KIuHVKQmK50PCcr0jWWgaIcegcjE8Hx/x6+1bpDGQZXc
FQUHiJIG2tGUfC5US29JslCFrdGNK+dzZwV0vFnbtP4//l3YqTpUmr6KLaywWVI8
7oISTTuldhqPxv/icZkO6wfniPWjxkGTj9YxTqt2m8/2hjsql664oJ1Y4yPNC64U
7QnGqKYETtbkPnOKGtnI8rbjhu0MAdcVm4kcO85CcpFtF+VKVSHJcPPI4s9DOW/8
/St68j/OIKh1Wdcg9i95RuH8KA6rgnZjFlGhfV2QGZEkYIvz9Ybe7sLSRBNQNG8Y
zCYxvfnxHiiBntYG4LCe/5Wo4cSCSCqASCzEshCtjtM1sIrPPCp8pyun1vzHfgpB
LQqoXVxA1cahm22/yc1rpDsTX8WRJqjUZb8lgHPfFeoJKsmB87YgruFsDKn8uz/r
LOOUQMJxYsobKwYu+5IPV6cZax/d6L42f7hPEnCUt2o3JdO70wfp/nGaCVWkex9N
rnZ3+l5bK0U4HVydMIOXKkAm/cPAT3XJy9xXtp0pm9JYVO12HJ9U9P2gMqMNF1M7
gPLcjDDW/6aXw7//zndKyD/PbDvfxyAr7aEncXQ2cQ4wZqN2BlnIFWg8IjuvmTXq
HugnO3gn5VQgXLHRufnhLsfxs+/RYMUMf9dcKC2KlIOM+eQPeAEoV1SbV0jY/sww
Te+iXejkZDKWprb9fO/zB8w8bQLBrZKAKGZUao9NdiYFT78B4ggkSB+MC9ufHyEY
6/mQMbNZWXXYijP2NLbc43PvYp9DldPHSIWqlHPLji041DFt7V9ggIzaaz/MuXG+
y6WB2HedrLp6xxnbLdLpaflikFAu96qPJS9dXka+R2gzqdRfRNQq18hI04eXGmy9
jkYUQ+hI42/b7i+LL7iN+fi35ZC7ftNQySUfdVpyIxi7xdAsMiaIFJrfzEnjkStk
hB9JL2FsfZCfAc8oAhmT4wcXIso/zd6PRdwfgF7A1OfRqSXb011wXKIDDc0Swqfh
pPzNJWcK97gtGQkKpC6RewlpHyxd8bblfeKD4rvZ3fqM4QsU93f8ydjPmf2fCQ33
D/0OG+p/E4EACi84/6Q34YT+kY9l/jip2TYW44uBb4XmS8SMKoucl/cZfNwUvZcG
1j085hUkvBYFX19bWOSFzNsjlIRkybtsaSAciGdvyK7qMpILhvPGAiCKWPa7xIdZ
ilAJ8EM3GhjOcyMiSs4wzfnSUcC6BcPSbtRIq38x00CJi+u26jvoqcqlZp/uNwlT
vQEWF+RgX1OiyLJB9fq3EFeHrfCv9ivk5oliim9wSVryW0qs+ABbTFXUv5IiIyvA
ZL0mVtK7Sy/TS9I8LHfvXpEV7s75zCEjYSU/VttmgtVEwv3YoedcdE9kPX9NWs0n
iPKVk5BNwJY0ae6sp05jt1qOQec5TyuWNUl8v7ffQ1Mb3CFpXvXsHY6zoHgjvAQc
Ck0U/pAXGnV7ika57LsP7U22TjopBHQOuVE5bWQqPkSdvAs+PmbLGq9Wm1vX9Qkg
73ZOD4IJj60gWmQY6hSVjytiJNAwmVrZHerKmlRYP4VhER9DXjvx4B8gW2GmIH4h
/fgbVRv2o8f4RTapxm89v4Cu73DlwUSzGxuDYm9tLdmYzZNR2KVqkc+KAUQkb233
kEMt4Hg6uAis7q2Q2JPHrj2Xtsw+2gNxiUJ/V1/QGO7YkxmU7/Kepi8r1Qjh32RR
PDr73KZ/9LqlDLCIHe8BW9ZRspArtf/AYsQbU/UL8eSgoJ9wLvJ1uHuMp3skZIHZ
Su3FLZLgf+P4/EfSiO81ifnT10wdWacFkhQhZLJa+NVSOAWKkMUc+NxhuHZLIiz/
10YRHBs3Nd6LLo7pChDfcCxBL3NWUtZFV1QE4sBAtEGOdFsDcTOD6uSKKXFaczNL
nQJo5IaT6N/xK4lhIxZXsF4zE7GnFudRjbiTOW9yh8Bvvjoj47t7Gq6YBi6ETEFy
uWIiNCL8fyVd+57TEkEhncTlgWiOq7W+6cBl3dYBFeZ+q0ntOeoLyDAJz8B+QRWO
bFQSd5B+uFzLfsj3stDnVGSR+2B6l5cpQ5Y/DRyTWkpzqaXR7dbcLzQ4+sXs51iF
Zp8TEphn0qHObuTrKY0QMyVzbGqY5NhuKXzKGyojAxlYYwC12Zqp5h8QNwHoQbS8
Y20bt7cnuzKxqzyw/OqLQFNJdqutAO4xy8QDX6H7G6yeLAjLQvbvI2QxHS7aXIMj
OXp9ZLi0fdqAAIW7A48g5AoibSY0d1lM8OHaD06W+20KlPgqTe6UEYREWbWIIhYw
JFq9GC1i8vLtgJ03VdpLk/K+hwSHwSMGYCYo2cXiqVYg/+rY7YHkNV9NHH6L/VtP
mt1hNFk0ythxubVcShOS0BMZhBE7HpVZodZXd/9wbfOQocswBj6EpMcQLxGhuOIf
VOlQMjkL2KVuZNQtonHpE9JEbmz/gCU8Am9Dj5FW2H2qUJQjcLUEMsDaP6XPD1vV
DHy2P59QE7elrlsj1iVS4TiTJ1EjmsrWSuubPHLVFCI7UN5QCYN2sZQ+kf6fW79r
jDQHSyjrBq4vqEC40Hi8NgN6AVwAIL3BDkfuCbscYn445Qnz+RrIehh5rDge97Oi
hDmPoru2akSCjWzmyYRrgmVjAhGKb6MTRYYE68mrymNQQAfucRGjKejtTfagMVcP
TWPVMPCnGIrhqwk/6RSKxU9i46g2K0zt4BCfLx0B5QJVDWMOkkHaayBTL9TqIyin
CkrHJmGgN53R1Z5h6dkrApX8HXa9S3K2Mf+yiZVEeJ8iNag3NrmhrCSKycHSIbP4
gyp2wnpsE7LbjXuQuoWRYVIkPMegjRk934pC3FrFWxDQogYAznGOMPcnUTu1KEN4
gh6iyGgk9rEUWTprZziiFHDOYfZACAoO/iSXETMla0FnwHv3WmyZcbAwCV3wnkHV
kkVPJXyIH9AZupAWP/04MZnYQsXzM0IKMBvAN6m7BLjxDk8WQTAUsG+zTfVsv34O
sCemt3nfySmQSQf8EakI2ZInFdcmyznk4AT3M3T7++nbaoBJoeS/pDUjN6BBkai+
IV34YumS1PSBBUvWE6CdJFTmGw/w5WbUXfj4s2rNXkhcZmxi1LX+03UXzxrIbr03
WfYKyrIj89Pa8fDl46SNb28nXN+CBO44jX4/eLp++j3ao3q6kbPSaE24XuzXQJ08
Ie6Q804KLrJg0vgjI6OCHKF7vPFeIX/UXFvmgDVqT/c+c1m669fWrVkPPCGCRn19
VnHWOfbeyYtRa7TUd6bZPGAmsDvf6Lh1I/KXmd6HVSvIRMgEpinZIwT/lNrToAYr
7sOyjGK9FjKgc9ulHNXERDAZIopH6nNULjmRHlnje/gdP74fY7lBxAErvpaNNL1y
SEQauz3KjasQEXKe/BdMHPF2IJiB6jW2TT1K7GlyUzVhsneXmDLS2pTZO+XI4haS
MJ50E3QvG+nkCxV/Ei5AZO69qI3pwyi6Oo83IUu610NiJ02y00WRA3r2xRbWICWA
2Q3Q7YeN6JnupJZrxxkRcZpSxNVg5crsDFHOWrcQ0lWbhCugb/ejrC8IKuClIuGL
Gep5eZweh2c6siH1TuHON/m48JYhlfw0HYLq+xwMQb6vPB13k5TiZXuXdnJYcURM
+ADupOoCAMOzBA+O2StKnivg3DgJAHE4il6u00/LnM1SJj39lY6ojQO7w9Jff/SJ
AIjq8DFxgcVr96yV3Ik5aec2wZMp2AEdSnVftwOJ1CZ86sD9JEALorc69O/SMJ7t
nsy5WTB4AO43dkxieC15To9qSrlHEVeWM9FbfeRVm4pPYGhxh7iSLGLOZ4DIwk0o
r2z7jQitzDie6t5OtC6y6wBrKyPecM++SNgSI0MvBkoHBhdnuhSRfJ+wLkoOpO1d
3Yoe2HxUgDEzOFEQp90X1gxHIudl9LS0d5AWWqcBsRYbTUfmsfcyt1J0q2m2EaAc
TskcKjoiZC79hZnRtTJWqScCyQM41jKeHS2SdYbGWbttMB/vLgZF9pWf8BOSZhIe
JWxk8NRK91O1dRv7/d+3LeezlRmH7jaXzvslmX3Ys+aLy6diUc97yDuUUOWeAPK/
re+qyDyA1hw4NlHPazxj1uG/G/9y4CnBzEQE7TKjTLOgFxoz+DB3ALD3gyiPdVkp
NbItZOx1kevn0RY0cjBBnwjU0vS5Vcd1rxvELWQQZyv7ExPfm0iIoJ4hKI5Tp9JB
tmpWC0rnrbPk8ljmuy0FUHxhBH6Q8TPmVpZ45xw3csDm0gOZtEcB3fs46GI9lHPz
HJujoe72OxpSd9Dn2niNCW9S9GbN4qLZFpKKtXLsP3eMPpkifNHee/l90HsWLMYS
T7OUr5f3W0CME/ImhQOB3RknpRFJ3gHAdQr27stvYY5+3yT6utxlwPdefc8GPnEe
hn9gROx29ZgZh7aFSw+KGiz7CnTb2mnO++eeRo8Tf64X/tzfxwJcZpfMgfuqoA5B
azMhS1/tJ+GWPnEaURO63jkAkzsBoG/jQA4pg+1Nfr8Zu2EPVsbiHu0+dwvMaHbL
8Z7ArNLKl/FM/3zKNTnZGegQmaXQTvV7Dw+MFMPqdCRqq6N4r9aoGckgdrSOKnul
TgGT6HaD6ujpErBF4NYec33ynpIs/S9PJKgQ5kKafom32865Tp/iC3bRoWlcrnxE
T+2N8LMDiRT7YmmuP0LLOgXyTiQy3qHHvxAGDZGE7HCvlwvuJ4U8wq8h8S6oL1Ca
vzeTdRBaOIOfDrV/LFR2DhHy6Thn/pTtx+d4oDd+pMF6ZGdGaNkJ7gP7zeQ2XoxZ
pZWRm6rkwVAU5itG7wkzvwGXsPL0vYTAdzeR+KUxjOJZKUdBNDwAGH4P2/i4dUqi
90JJrvu1ibr2IJigN/wa+BYQzsJL4bpXTv7xQ8I8mxIwPhSKN3WJlBYWbqPXCWpS
R6z6pRCGZn9mmKMx+exTPjDO6Yo5OzyvO3HY4TZHWhbogTyXaUfZ254ahPQuyWZg
lnToL11pJ21iZ1beFKDe38gmnmkYcVUYUBK2HlUQpfQSupQJU035r2WUhSCyLO/5
B7Q9XDnBSBWDcSJkdo3xfL2tzPTmOLgfQ00UNWVkfMjWwO5tkddO6RslrSxDlWg0
X8yCYuMQrM/DQsdb84aNeR8SlAulAxLL9q0BLR65qTdn/xjErC3pqKqsYyBibxwl
Y/RxgKKW3jS+Zniefh50nYxnosKiV1hklfTQlL/5KYH6CJNI6vD9olEy+WFvxX6V
sdysksjzYBA1Vkyvuar57yKy+zlkTHXcyEiFzyG0GOPwKqGkYSBcc9QB4du6CYHX
mMszdnuXN96gShUL4RdboI9sKH5o7VLyz0cOi70uJUA7p/KF1/4HU/yx/NgXOcLz
f/LILlTxuyb5tATfk7NTKaEx3HQOf4tBeiulLde6dcWs0kcWvcIHmBH48gYU2rJR
tV2i2LcBfoQSdi2T92ZAMo5hDp6hgt5x6dDZ0SXLdS821sCgkMK1yctDuyrb/BXt
AwqlVfRrSEoCUYHxWK9282ybEOadnmcb3ZkQGBnQ08DaPU2ESfHOMeE2jH427kka
EWDAwyB0ugDAZ170M0SUeQAUs+c/pYzH2/NXnRTYc/YH9S8FuP/4YSVfReYp5Xis
z/k/Xi1OAIjQCM5dmyr9DrT/P065soC+bFfS6grKY4u4YOR1+2vhVtYEmOnIgCm9
9XoIxGQrAp/mqT9GOY5rwOOWyA5IJmqSJw78biiakY8CLaC9gK6DEQYeo3m3a8py
Rzn5bWy5+JpAv4pop7Dsyh7IXrNGo0lvM9bYdJJSBiGpZpjh/Vz+sl9G9cRB0O9a
oiFXc+2IBMTlO4nhH7316xYkzx1DDqxFG2cpUGX8BMIYdkpKqOvZavvMMJESt5+Z
bS7NTVpZRvm4lcUcUr+oPIhj999GTYsvE5DwrBKvxcpxOP3yXsOulMLmyKgsrjaa
9CIt6RsS9b8yLEZXb50LnNNVcA2Y7gWSvENmoLmJ+7WP3bkElZ7W5d+LPwMEL9Fb
M34KWYIoi+6i45xHwwpus81OdDnDk9Ny3f4Q9rgP/fwn3CFdFYy5NNlOQxGhJzqW
bbjzjwHXBS5ZBGWuV7VMxVwhvrmIhb8jmJbC7elZZnnPpOkxxltXuhue6li0X4My
UYpS3f9EL0/JDtW62E+mtzlWgEePD9c1GG+f9ztZf+8G0uSY5FbKyOPYVZlNxBYu
7bcLzjOliyQB+03LG19JclRqc2tH/yo8A/vBLnyYLGeugPBGlD4w/EnR/qJDiO4l
L0KTyi8WFPDpFZCsjqSBE8LA9hnysYZB1df4ZihCU1/cX6XD9DB10ZuWwXQwIXUg
aPFMSGA62aVe49P0sC3bk+l7kS3mr6XZaNVterAhe96zIJF1pthTPpmqi2SFe+Bi
NVBlNBdgw8lioxxHfyaAn1qDk0EJFbGUE2HT1dAOU2wyqBfa6X/FnnYxcdbqp1Px
mqcgA4T90xau2UMa562Rtiq48s8kqQw4ekRyDTTOHRQ2kGdlsN0Uua/yz8ZZv1d0
hczL0AkNJOU2IvLRfO4NmplEVL3grUnzOaMTYckqfiCufX0Y2X3CVLEWxAkxNJxt
3HYgiip4pjixYPWZKQROjr9eV1X35oYnG4RqwZJ3tJgafqmXvgkbPqmfl/fT7q+/
QfgKP2QjkZEDit8d+tzWcZN0tvp7bksuwNcP5APgi9VVN/H5LBNYM5Ao/4pyUts4
duyqXu0QWAPxh69Ue2uHaHbCYVJLau8x47hafQFwgaWOQ1ydmyjpL3aDnF+E8pRT
F4fN7lhpK4NdmDyC7uwxIHL/DeH+3G9124x6aGOz4rXtSlXAh7hDTD4cN9rlI2bp
fSm/BUdzmbcVe7BuzoNxWzELlfoR6fgV5BAU0R3sd9/+W68oaikC61nZzgMEYn45
vEznIk64Xt5GUpahwUZQcB/OyymBkPsQi+fUnh1omEu9RiZ27uafuJILgYhYUWBy
roeGpoxm+8xWREsie8aYMMDxuvQUXNv48XUF7ECCz/TOptvZvu0K8GzrNZebP9hB
3zcw2b1gHJlZwMzfSsxJ326dh+OiQ1tIEhIhhjfgiHC2uz6EsTytYgl7hPCRnIp+
xw0GbD8HBI8HoeJGlUclwhphddKOmTkql2mstFt2i9Z4PPYYgXo8W/yeC6iI19p9
R9HFAQ30SmJqCLFOLJWEB5l4q070OIti9cu4s88n7XMQkbUlYZPPNsc0pNCvvar8
rA8ID9CfQOzpY3mACJDjOQdEjNrkSDXYCSoM0nVOPSrNWqi04UqRRt5k76l1t0wB
G9ccWQ91KiCImCW6pQV6LraOTj+XEB3EryOka31xjijZikWz3gV3w5Wfb2gKdkJ3
BQpOKv18O26f7l95FQkh+1PWYv78sDumeDbh7FYB/ptKfoXo7Lb/WGyWFfkkkobt
JfDN09Yinjq/yC8iP+weZ5hDnqoYOGL0ZZKDdg6cSVAWF+0mxuGqXonkud7xb5MW
HaPehTIreV5NH1Q+yPeGfFAwcYXmixmbMl+Gf4TjNy74/Ntljdb+jxfsniO7Gccm
qcaLvPSycwub2SfWK/RSCRfrr2JOHMftWhWMgsI9hK07y9ym5oSG9rOMypCCFh2H
ekRVjAiOB8YJlysNhxoQLMyNAqy7KMI2wpZd0bnMG05v5jia4aC5CgcdqwEzRdvr
8E7BCfBlSi5jB6P4PVZmlSLQrJqSFl+G7k11qK3J0+go19pe+sdMN8G2tbU6l2la
4ZiYmLvz80vBg9q7nocZYDhXQul3S698vzD67Q0Yz3K++W5EYdAVpRABRE6bklGi
BZhy5yd6ynN3Z1v8PnPcf4hFfc4JK91PS6RURIy6JXXvQbnGGs8VKEceIBKK5kdk
laqz7OcXu4hAuq/K8OXdJpW8OJ9elQohfiMkKhCicqJAL8DVKZ8s74GHA4e1kQyA
+IBs+3vdy4dpn+jK8j4H+08rI9d/RPEYa2lTZMmrzxt9MRlzmH5UIVMffovEhLs3
LVA1iSSUPO7/6/d1C0J8SG/QFFjj3DWPggKfHOtUTBY8zrwSSq2CHM/MFgqsq/ke
NBU/kGJwf7k6Pe+C6u5XuYrcRbWWcO8C/iuRAau8dBOPwPReIFfCL7vE8a1gVEhS
KKmWW9+IJMADwss5GY+fxeK6aGUJN0YX7QtvEn0GgcOsEIJEQPoxDvOHePkzgeDS
/QnoRoPIF/xvgVqc5XoxPhiUnJYOEIgpwScydeyP3c9yzia0qb2HzOe9KTc2bE6E
PZfK82KRjC0cTrF4a8AVVz4/7RhrmCm0vwv2MGZ0kUo9qH5IThjbuOM+dNtvaXVq
6v4BdNnWcssPyKr1v+x+Sqg1ZAS1RLLDlm5byxb7ZQixmw7GEEQ1Be59984/JM7h
/hpYlGEnSuUiRr3pDQqISpHL/Q99BprHRTaCbKHv7iCqhCeU/Xk0WwVycIh8izlM
hI7LXk2llFQOtgFjuIdVq3YO1SrK3ufIqS6XxV3/BKrAnHkY6DBlOm2FUruVhnKq
W/NbX1PZ5b1EPpKkDgXOkhJtiv1eH0aMYkrk6fK+HfD65An9ZwxAdPLXGGrpCQ96
Q6ffiVsei9CQ/NKXXyV1DavtBY51dpzCA+pl0hmHzxY+ZDOr8pvX6gTpbUM6Kpfe
yxi88XstfITGb9rEpOglL+i+Z0m4A7O1XFYFqAc1dSYfjb7/vqTYQyWv7J1shJHR
0SU5yLWyBxzN2ucRNrUnM1/AeP+wTpBabcsKAUA1c8DnJdeprhF6Z164n/UpGPR5
4e3p0Umg/mA2YRL2xE5L0hFh0lSMh2//B+3KIqL29y4zY7hnWcxALOJkryNf2wNP
YzUnXmznP/SidTc88jAP/6XC9KhwM14hHT8SNexkXJ4jOjJmgAanaDtdtr9PZLu0
hyyLQepPv9cKecNI5SrBPns+YQBOngQuQ8pNEk5REYD6BiIlptAWt3wC9zlMhjxC
MYGSlyhoRTFg2QAqZ2ztYaOCMUecAWhq0DSj+vDIMobLMWHSD7I9Tu/S7wLkYkCr
gNE2j685XzyDtEW+kKyBStElvR47HdcuyOZjR8E89B3LdqbPeB3OGV5z2xj1wqeI
rbD8xW470XTUAwv76ilatSuvGMcgg+fwKVitWv7rmOZAonarGsIWXTCBOraIb0Xb
zOJ5x9u1ZU1nPqw5weItCHzL44RnsERP5JazPbz2ZEGTzFrLEKtc8ocFSFxmR2Vr
LPcwWoY8gB6shIB+iz9jrlICAIHr9kbyPEvJwepCNkKIxyoj5pJaEzARzoXkQGFR
dnPvPcaH4dljTBBu63gYtDsg10zNfVY838IbcUpS45FhOSb6bww4hay+yVUfKUsx
vi9WCcU9Di7DhEmRb2KwmwjA+CmvIqL+Zcf+qA4oV0kwCjmR7grSMBu53iE2UCXr
rHo1XHoSQaF9cSWcBIoQfkW68W3W7/BFKGbs8iAdfbk9GrLoBapaK3UXDjWbacDe
c8JYCMZ2z7pRpsJ+4DeMaG6D8WOW4Pq04891FYOrIoYKlf3yswQxOx3RNb3Z0RW/
bYCZOGN+nGcdh/l6JQeS3G1ogcS1XGWC2//V+5CDa4VXs+OlreYNqZ+Nh3M+tir+
0lUtjSy5kokte1IMnFlFTCSLvfdAOendccTyheV4bUrO7ssN/PWz/ioPLBgIuEHr
h9gBJs4I2T7yU7aIEB6v5mLjaUVcRbmuzj84axirh7Hr2DTnsfy9gOOsn1+0Swoj
GRWUgIpjYCEHW6gxkUNhQ8kqFekdRr0DhEI+0UHAeseZWcJ7mhgqlIahB4OxbBF7
vrgDARxPyf1+kLrOsLZ2TuFB4MPl15dvylGlPBm2lqmrFWwjStxx4fdsfsy+TUd3
WU2vRKjbB0Y4SgdERY/S7wcHnT2hFo5ll3BOQn8tBY/PV9xrVBiwBQGF0+W2lzCh
adWuUs/0zjJStOl+VTyknJtY3hckuN5yEs6k5XWWk/SCFmi8y2YMlD+5sGUN3Phx
smnzKD2qwHkOdMUMzmDjWVITWrXa06QpwkXnKA4cgMQcZ81CgFWIrRHuieKLkayq
z0n/+NJS+xeSrC/dx0GEf5Sph+TAhJjJ37JcE8hZTyawRTanzK7SGNbZdC3UMkui
xPNps/ufcuabg7cyJaJjLt4xRdZseYdvTzLtALskSQFGoX9jit+CVTwvDJbMI5Eg
DiCy6N/6DxMOojZEXMJn/6E+FRCV2+Su5t9PJrgC8CrP7KWoWgcnX2HRU3Pbd2k0
R/Im0xSbVWXE6RTl6OROIHvi6gb9Q7bbhT+nfMIQnDf+kVnaE0jF8D3lU1EPF8Z8
t1JYQWMy39VG6QmAkayz5pDIsdvawRSQC0FLt6FaOEEdZDbQr9X7Gdyt7xB3ayyi
3IfBgKu5KyP4jIwIhcIBgxNoN4UO8o5p1/9O6qeAtb4VQeTa96QFMLR/bhqenUrP
ZY3f1AtwIbaNBWkMJPsRLqfiAaaPio15nsdA4WYFnWctyAo7HVsSMg1ZtCndVvEh
f//Ew96MVTwJ/Xd/3QpVy6mKOf5mo9IAqd8qPx3GBbkobt92GqERtCoDmq6MH7w2
zvW4fcVK6YV/fnbITxw4g/2+JBaF/dvBC5VJ321ABwLs1S9x7seymk+zUi28J3xO
XJ29B+S+xtwjihoyVql5kSaWbpR0NxzpuTzrKoWTmZYs+K5Adu/zr5XULVT5Zrwn
LWRdnC0WKPzhT2c0nseVZuE6eh/UF8qY8IgV1Wnuw1MFlFIeJEv7zBYb2XfwO/qp
OIJJoFjgrOqlQrcAZ/NPesyVWAsZ8iw2SXAKRhnFV3TRl7OYGG09bd1OfrZUPWqD
bQAkRi2S+5nbt3bbBc/T+Oa/Gq5l85JxaBhuJD8GoG6IHtsaQ31J3PXQKYPCKrVU
jQsSpA0w+QvAgo4FCsChxPuwmMShwSot1dmWxum6f27ddH4B0+3Y6D3XRSOg65xq
PKWhGKeedzhJBJJEXqdKGdXNkhlVf0xBwr0nEJy0Yr+vFZaekiw0T2csQ3f69oWd
mP6eYpoT+zbQDbjgPpuHccpJI1A7vqhRTMdbevBXLdkGR+PQW660DxWiT92URDxr
CFEzW5FZnDfjdXxMO72nlw113cBskg9qkCKJ+PpV8CQGrOWsOn+JWexlA3fLc94n
Z9WF5aTv6iEokwWAalBrtpveMQhBap06jH07YPRy24XuGQ68de4RTcBTNy4c7UpH
9fTWCm/NWtL7nYt3tXY5yGhwHMnfItckKogeGP9wp9y1YOT/eASbOoHMKFybmOyr
SyDw5dIRmqk82RaT7pCFsEZ1YVqYeJH5V7sM6OHXp/C2kSTElWk1zzoI7t9hdC+e
CyCKH7WbAuWibqgdREVbDFmyktCU9N7lU18kd/38sRqxMhmoyuYSB5tIEGYshSLg
XGa8EGGSv0W/2jP4sq1rLVkPXOdCcLDs8e668pJOVNo0BhKxv1aX6uOi7jOBotyC
fki/udvB9xAXhkDuQU/imQ6tI0sT6l8oyRh6WK9bNKziDYOJV/uf5STm+cGPf1Qe
64bgBCj0TOjXItfa8bt3/TARzfwl57dxhk+ow6hQMSdlPgwxXkayzz0jbF37KMRS
lUapnM0vBibRXoz4aelSSDoWi5UI29NEppJA7fEmiDPVcGzFY6g0UY4KEj8UWgID
RpfgTxQZfaZT0WWfluvWrYuYpzyn/Z8iBMTvyZuEqhsUPTCJBFlmtJ9x3ZeksGOj
SWzNd6Zm6jP/91doI2DNxAikiQah8ADfl/L0ueELrIyjnxPwfMPKrbAZpFW/g8l2
AryRMZoxTT6FtJi7o0xNHPA9SSvC7R6AEwaqe3glZObWHVB4QbxeOAZvq1MbOBlp
gxi9FpK46+5E+SCl1ywcp5K2LoDcuOi8c5XefpU751sp6PK2jy25VCaHSrj9xWBy
F8eLGYCPTEIkmwpPzUtZ6Q1+mNPdbuUwu+D9SN0U9ddlR/IW+jqKs0HTSFHrbyS4
PhzpP6aB+PlZedEtc3RC3v5GwiVtwIvJVIHwdst4Dpr2s21/ee8cR+OSbSdqgX+e
iwI7qHUpQ8IiVHP7Fr7WguioL1h7kb1WqsYZLjaiSrsDStMSl6I4cWBmoDeHjamC
WENwiaG7UXDMAe3NSX5E5Divz5XvP9DebwHwyQxsqK+h47S43tPkfmZKS/h1IrKa
6aaCkPkhmdl4Nx4qH6Wbwik690Tfr4fqxxgPyQmGd9YgPBmOTr4/kdXHQQClhLGi
iy9ySzNJHfo0MbZaJuMrZGqPrKWLdaNmehOB/Y18mceatQMeS8r/5zu/krDFedLK
yZKXK3s3E3oxfJ9xVdyOHaOKCrQC0y321E1PU6ze1VLNJzQ/6ambJGdpvsz1fbnU
n5pLGpRIJ6oiaMU5VJCqYlBC9QMBlzEcxJwO5kIJW6UjfPyfQQS+9dWcoSxeAxc6
bPQZg/Z8tFFdgPOruoCLhwy7XN6XVx7Jhg3hO9RM2O0h5/ahXXtTSHlbIWVYR5xN
i6lWl7wqCN3WjYRN3wn/FOHBRR69ccXeos7OspV+jdNy1rjuIm4MImDxZlSYEPuK
5oTgDdG/M0sn12GL7kcoNlFL8S9MnPei0wKc+e/aPTwgQcQp//ml6zT+Y5BQgHkd
GRKnfsrPJ8lN+PNHLaxc+IWKkd1Dj6bP2MFdaejuRoWyCPm35uBTyp5nP2sD4TBS
aCwC9BNh8QeusFHTwzEfMP9YnabVJ3BxfodxRM+qRd/6fWjl50XGVEcBPpd+S8/t
6rHb0cTWrfTAj/+jsmZiqAODdhIyjdNewxPlolmZprzNxAs28lnkcv7tH6Ii+0Tv
RJC8RNK6T+BIv2ZWU8uv7yTS+hyqIR1edjISTFwRZRaIHDbAFB3ajMyD9Agqjwe+
4OQE9cGcVVxWcrQq8WQ2P3IKhLDb5ChXNAVLMFQ/Tn3JSNwjU8yc0lIMv9zYKkyx
UyC1SPK0kNO8CfiG5U3qC3T0Xol4c2xiKm75x9AszKDTLfgSiXSSuKbQH8bbwsNk
eclr8e4F2I9DdXcVNWueY9RZTFjNA+++lknw9a0BA959S4UD5uH6527GB08grOuf
l4vnDC5xfsmvLYH3wjV8/Ey0PZxWxJ5mbvSy579BowcRh8rRGLMXD27xCbqSXuwm
4AmGngNnrAPFmBvqPv9pruOrOfJdxjspegya3TWVJHUDnHd9cyrRnXj1MQcFLZfl
Hv/u3a0OOJQPoHyPLDaZ5cTeIwh3C4nBwbCVYexTvEgQXMYGhSmgLTueQGRfOxNY
kOFh+7ZD4ji7oKvNZJKgdVEkEQNSjdkJYgrZFUCzPbJsIEIJMzO+9tzBUNnn3d45
g1eCaBfY0I0Xmun9opIvPCFlbiAnv1UE2fS/oq+rOs2Fvc8c+flrpDVJ+kvfhw6w
L47sSDFFfolGri9Ae+pK+vV7YUWVDP+6JpKzDD30d/wGS54IDY37L7glbk6alu2t
paLPzy3eNsWBJoYNQGdt/kiYe9+JyBBRfndyRSXiohuwTcqBpp4kpE+mMmSxWlB/
AE27+cJpaTSEG3WX4fps67abI+odFTKbk3GS+maK45Mjq2dMcZj24YiGY2CQsleh
RSdv4nVt4wGK7S0RKJHire/NbcI0/Gh0V0N+o3ra2mMct+IlIULX1fzHShobFb61
EiNx7q249cdRF91BYC7+fFRAgpybgmiab5LkvuUkmeyauqUCNjUPRMsrD9auCcHj
VqwvOTXETKNkzIu/c7L2g4rNdB+LsWpsBjDLrSPbrRITqByaQDiFdU/ppqu1Gm9q
GAKKY4uCTuDNNKpf9UyAc5T4MwTUeYtJqxDnm9XQlBBPw8HaYzkZNTRdnTtv4fde
1iYLuFiNXBNGKhlbSqO7E/MjKbJr9WR1uwq7yNJI07o2O8vu1/puPYstYTNNEHxj
Dcf+fR+bQeIfFGBZbkFFO43rPzNsaqTMvmYE3v0rEOBcuse9eCVVwF3hORVVnoAz
U7A9Ksy7dlU8vwzekt886CEFb2kRz5J90xmzaaKBzMfPjkBL2cPcpihGwKrdfmHv
r1qC+7YYakz/IIvMXKCg+hK8HwHXuZrcbiB/Rco1/9NIREvJDqcoWryUToYIYsQd
H41BSdqLHsvV5CK0b6OrJ0oRxw3YVczTan8j5z6uyqJgj5ZwDb1AHiJlk6NhC1m6
bk7JIrtgaUrFUeHgZTl6YWRg8hFBveUiLVqUA84mDMiY4s7giTgYjPV9f5RzCRWG
th5T2rsOdng4+mEkCx+F74C8c+/dr+9GEO7ubcTEJKAcn1nWU2mtNHaAecI/dYAC
0wXtvYNOCrzN5y7rMYrK6pr+jGxIkzQk9aajj+c+lBU5GQqizRPP6oEmilnnXO5g
fW+AHuLpFH7yC6t7TlqsIr9ezPCjgR5VflE9HVj+R1v5IbCCp8kj8iv+mHpmGfa5
JEIINFWq37JCjCEcbNXrAgGDs1ekNQWcmgTnQ0lA5qJMfAnQ/W2lQmEft/b3zFYv
d/LmW8pnAbBLhdLDXMKHHhRPDtUDIr3/XgPOOemfuxpyk0uIYClWQOLxec30GrNG
SeGxUdUesUb0O9Y6KUeJVnMl+vaUav/GRh5ANgXnNivI/yIDkguu7JAk0undRQzs
DRuC02kNRyyShwRy6AuZcF2wbah+E+6Jj3oytZtB+HhCoxUWTOHQbADmFPEPdVcO
JvEL+T98dbz+qiaVfr13HSve6/nsZ7NuLFoRU/2+cnBSY6vuZPisjIzCiq2o9zAH
F4YP2LXgUZ+ni35qJFg+8K0szwLOVQbDa7Ehiw+GLocP6tQX6NDkHUPwiPj66/ps
0S5HMcO1IsqK3DoqaFlT2pakoEy2eRLgVLJqZ4OAWS+DPcsUr3IZOhQmt5gqZxSh
LbZdeUrPVwZaRwWJn2uNC5y5IJPK0gdjM2yYnTECs6EKxe3nh7U2qgwBN1Ce5xZ+
eecUPaawyISjwa8SJzLsGlt9hBhoitckU/YgkeOplkDD8KmDw8ss4OzIkltFMeRx
PKkdfm9QQ8do4wfp2gImYDu9gwa294tgUZvOOQDT1xVbw79DQZf7owexBR4r/43B
lI8sKVUVHzEFTnXf2SSC1NhzGsQnJkLjy/O/oRRu2uwux/XbG0X5xMAMTLL3Ai/z
/zXvLOBN5RuK6u21CjOVE5ukNFtZ9q37bB6EkkS8g0zhx99zjb83ITdUDR7+E+XZ
Y5fCroukFPycKIQznc8miHDEqwLo6kEzGAQ8jPfMNB4M/DFjhJKQiqU3xyGM5Zm0
ZKnyIQPXhDMhsO2JQFQ6mQNVqY0dL4qbd6ysZDpqVTUmJBQcgJ1EcEv9UoswgB7+
aWaAFf7mu8NNrmbuotohdtHYDelbzR0EBj3RBcwPiWSngO7DcT1249BlNN5latUG
pHtevT6slJo7GZ6/GGXz0k+VWouJxKTCH+xKTXOVlSjNJotJfUOsQ/VPVchZuX2j
QFizk10ypEQ/hmy7YgusKIMyMzrlyzppZ0qmqARIAjQrMnVdKmwdNXLvVmquEXEU
naIP+a1DC+yLKTS8YtC7seLTPrTa1HXUuofs2b1t4QiF9v8gJ2bPbodrnBVNgig1
U45euDLVK76eR+jUhsA9PTsXGfPHXwC3jxnfg5N60RUtxihBLy1LvoifgH2aHxkS
apgVsrCztn9VhjAvuS2MnWTH3+XalPUKDrj0xvw8fL2/WPsnx7kx6uUxRivs8Di0
MUlMEPME8KC1zgzQF/04ldRTBbjoCJo9nH4FWHWtew8SInEekUU6/erlMwNNbQQg
LLmXrU45RZU2XSudDbcI/iVREvD7sYMOpzhPrLrltN5eesSwZoINWrVvZsLafBDQ
Aigim61h76xxzPvK7GwpiLFumblhfJViX+gvD9Tt7a8lNQHQL1excYY4mxNhxn8N
Sw+seTPDDh2CCAEB9tPrSrw16DLR6zXCa8IHoNLssz67+Q/2xPmGZFnLIhfCBwg+
wT9t4TStlSqkYCTLvYH4OeBxL2jxYmOjqO1RFqkIx7rJDo6Yec3Yp3prFbw0XBJc
Zb84Lp7OZL+C/sjiPK+LRnwvk1CoJlech785zvbTkEImjHSvIHwbMGYnKCtgpPCC
o8KNqb71f/FCFn04YHJjlf5U8VdcQKakoGIExTbUsXXWBOj5H7ZJz3r2rbMZCJMT
Xu6NqLlzaW930m509FJuHmHTDE+VyBLEA9GGRBWZMJ5AMLjfhmyQmmW6S6QfSob3
d25YjnnsYqEqhQv6Oo3U57pkKbxgJ4e43gx38ohoeRuFgn44tRePbNMKxJSVgVPq
iNp7jSF3b8ZEjw//Y6pAnchL3mVYswDSCtkrXfgJT3MaPiEf1atkHub6sxvnr+j9
8C1iYDKy7SM+b0GnkntT9uLIiioRXve/hhB3Bn8h7Vcq53gp0MdTPUk6vKmd8NpG
SG1HW+NkJ9TqKrTa4WkNZeDf3hwVBhfNifhWMzIzw4Z3JU+no3WiYtFFjTof+d4r
lhDEk22+2o2vu9W0dAkCmQw8ddkHvtYPmNPiS6/L5LOhLS1Dr1disPvgDnPa1ZCn
EZLFo9EpeNjePhRG47dY+KycLYXtnuJWzqoRwHuoV7EpWFpd/r2W/x7e5NKeMPNT
GRfLL13MuP52+LqR+/kjxZTD/MfOhiThAr2+qTbVdxe25UvqVMFOGYn8lLZl19OR
O4D3sZXWxS4l5eqBgT9IHSmKh1NgF2yNwfRQPkMpNzBEpdhSomo16YskM/vWA7yB
8HJBe5t6c/cGaujcMn9tQIfPw7MCS92epGAjE5xjfKpWXl5KqKU4DwAhrRx/d+X1
VtP/KkALppqFu7jdEOWrfUkFXKmhm+VeBKi3HdF7KEIuz8OoKFKm5zuFKElOAwBl
H16G8lbrBFgjkRjZSgfbivbC15whhZBpEVe54vS3NpCTQF0CTNNcnGnF1k1JGXBe
Nnz42ArFbUGPrGHAuzu3SwGPLEWRD/vIFpico+fzHbfflAXb90uFJW5zjF45WeY5
hDYIGQQR0QH91/HCZ1sIBsyrAHEQiZ2kKmo05dl7NdYPYVpn/APB+zVWTiUhlMpO
TeoClYxZw18PuGfraeS019oWeWZhNRag8O7HEckP5zAlXtAu7W8OCMtJafdwYolt
qD+DNcCI9UOf1RxrM9zt6OdCOJftomca2Sja5iJRrDU211psslsvYQvP5HsutNwx
3RiKQuPHWkcphXe6ZqdnOzke+g7ngc8o62Y4SLjYL67MlJZk6ipo+aeip1eZpoJF
XufmiEZZP5FxON2KDazSCdXqh1w5V8iGhfFuIgkDA888UC3p/sDvX/NQsoz3dfFL
JqkJH4ZPHpfMbKBgrNnZSEX2gJ1UqT8TXBl9gkVXIbjrvz973QDTrUTYpc9RBFWr
fzcSKdFp92mJqGgFWf22GWCPTBo29m3qHF88uI3UagqjdhH5gsuvR1zir7OgmAIy
SvfS0qWNazkL3jsjDgLOj/zAip5AfYU0pljTdneYrmuKcD0kbdXdc36O3JE2qEhj
bEBQxQCsk0+mi+Ly9HUINzSxOYVpdJA7yIz27jflG8F0m4T0GxrOlBsS5zaVXkz4
dsfoUoM4vXQUURmZd62ZTSDCNWlFNLCVTT+hrGSppCdOYHKjNpPyRr+huaRPY69S
hrMhf8VyenornMylRz+/uqOl2WFdxPYbbQM4JM16jV6yDrcjmNsGo3Mv2eKpX9vW
H0R768NAbV95af6Nyw/OTHqU2rqdJzYlHF3J28KEk9EWkbiA1z3Taem7YheoOWMP
Y9mQWPxoAFev9tHlMtGzbrMihgOE5z9DkR9gGztWIZNYAnrUXv/rFd/w7CaUuBXj
PdkvnKBJnUPLQbYLVCoH3EPUylGaMz2okFO7YsEgWH2yfSiSQvSIZcM4tkXkFS7k
gSXP63D+mfqIP/79upC5NHwyE4qr9cORtq7S5GIFdgSMMN33PrezoIBZX6t2CV9a
Q6cU9fH/7SVk9mp/Cyb0HCmcnc+z/gEmSb/aHnm+2ZOOjlTsRUwkC3WOFxyGL88V
ONFbGlqGB1bp5PoUqsLXnblvPmQGnXCIK/yVS0/uhrDlYlkgXabGTFNs77Zi14BI
rjtrX6d3JW4C+R8i79RhdYlOYJjmENHJm/nVtlRkS72V7llRl4iAjaPZyJHf2XBz
aWNgOKBP3DvoTwyUmtqoM+cUXh0kzoRFjkcrEEWwbE9eGRBArrVFzokck0qewrEh
/sFNKccfvs0IQg6YXJSazprgxUX+D8AyQL6plbOFzZMDTgtRc90zYBtK4aleTosw
AbPLYeNx50vwRANre9o34B8UkwN4MvKulhmXyIC1fvsgfhQEbuooRbTTqzVs9pIS
hGP91IFJvrn8bL5Ikq9UgvbewB3GFu7+AriLXcTCA1F+be30N5zBs9tqf2LxjNj6
CGQ0VV0X4pKbwu7Ws7NrS6SOjmkXntOB1cjBh/2FJypAg1Ogyj5A1iJZ/tKraxqX
5Pn7K+bPFM0AFda95WHBTYPE1iWPvkkLWtoZ804D2DoruJJSW1KUqf8P6FL3fOMv
vO5C2AYUj+xtXZICIROln4Q4FUnK8DiczMrsg00Glg3nAoflQB986wQsRXWFh/rK
N+fGkSXB0qHQT4BAxhr6fg87aGrerCr8lfcsZ7yRdNE/Dlnh8NjZV/j0g8YIjJMy
l5BTvBgU6+cRrSOdmOo1bWv0glx12J1HzVLCYGwu9LlCphGshxgP/I2V/0l9WOTs
N/Q9f1DfMxiXptYyVw+KzDk40WPfaQFaIph2UGyw86x0HdNFKdA0nkVg0EPd3rVd
V/h3V4rp1t97QKzS+okSiNXCfUXoInqQ5ba6doiRe6Rt/h37bzLh2mm7fFBnFt6E
9TiwWPtA2Pq9TjfbrnOhfJcKvEenPYofdorPiuXkI1tUwwyJZQ1zzAiqqikFvcQr
iUs1T66vkAQJ5WT721QE4tD3jHfpuJMniEXPL1gKFqmboY+NhE2vH/shjGuzjw9i
NI5WwpsMZl7UtHLPXDC7sFdPPdrjFKaOFMgN48Fj1K4syQgdbwyRVqaafYa4TP6o
3NpEfn8QDRY/rcjH5EJx3y5yYZvecfpL3k/cg0882w39bj3YoaMAAkq2EHNi9RL+
4q1i57q84CMCHbBPNffC89LLbqW3/iA02gD+HKFnVqyIOQWitYMzi78WVJ2fxarC
17uxF/zSRypC7l7YYIhfIv+MpCbbkw/9Ic6cT5HS00WtIPMQyibGnItn/y0LAGse
Afw5qwpq0LUPYVXpKlLWd+AcO8UjdHWX++t5PSBpctsn5Ek+dWo6CuPaewy44+XQ
OnBhEHg5DDGMCAo5LP/M4PlubM07KerrwF/jJEES1YDK/G6czVq3d9bkaQ4k3wPa
ae1FaNwjQigDG+RQ854qlOkB62BLo4/aqD3kEzfeV4FWd6vPXL5LnPyHnTbf8Hf1
RRd5+lYDi1C1SKROIun3jx3FdjTT5VL5UEtTR3TInuza7eXhZsEiXZLSyN4gwneF
FeXjjjOrdjklBfzL4qOC8hg39WLeAAkf6vqurJVP8hk2bGrlLhhnMPUdEVhBJNVT
rBZo04YCbmvJWoqwxeWtmkoyui83zXn6tW3jvZq/6ygcywTEAhKXREi19ltAzb1W
WNKiBd/fk3hkJFdutRcFQDdzYc813TSCxvlqbPRBOx5seJgW4P+AKnsUjvy54CqX
6Wf4uQMl47gmME1TV1atBA8TX3s8Ok7gYLVBljes6kDiYDdfoNwXFKGlUloNbXvL
HUFL/2jQ+yQxi5gmJ37xatt+7esFapnKbw9GNjfQ5IBogwyehhOmdEwKInSNu3Gz
BF1fOILT0Z7iAwGVfJmj4XtnM1E/r06EYRW9TGsQbqIYaIN6Pf2Mwc1qrRIE7AZx
EG8STDEwQWlysqLcK/9n4Qcsdd0M1gxoO2E3SFfw+6HrgTNPGKBnWh6RCyI3C4Ou
iNyYrSi8bxZNT2qUumpDv5Z/ESmBbvqshwqMCQMZACADVVYWo20JHZX4TmM2mVMh
8uCwJPjXXist1uFqLAvrCnlw5QN1hFZw5WVxXqWtlOK0CLwL+qiErfm2eobUx5Lu
vNm4oM0jf8eYWsBjS+B/bqwECG4/pbVNO7WSGGOxl6Av/QggxjzecDjkLnvccG5f
GizvwTiu5NG/cJP4GSvaciuc1M54V+XhIWAHDpxlXzjb+diOHB8pOwdRjifaR2+c
X8si9/FPKoMER083w+xiuq001Ext3EUBVC7mxadYFqwejUSfCoiI39j9m0gr4QKJ
NCC7UlCsQU1pO4iH8qkqLKLFSrORY9/HYqscFHVfcyMHdA/nXQTciu6Ccb5T3VWQ
6rMN7pxfQ243FoK0937rV/irb1WQx3Kf60V1kTrG/hXJEcvC5tZCOGmJGf07934K
P4NXOB7W0kZj446ilXZLjDE/BLBHdl7/s7BeyIa3R7FKoYwUuNC+g11ljS//jkJc
cSXsyZuShAL4nnHLkSvHbMSyAPdoGtjLeDcmsN3JIsPYOpbUwcIAfg+zIq+970VB
KdiAm3V0QLUwthaiY7meTHuO+cUtcb5mv355MWzOlL1edPgIM7S1KUp2fjwz0YWP
08WlKSQgtkMmSqbbJDbUxZtoAr/RxIMf4vq5slC4hw6aBDbvPpQvc0rmCqJNnPvP
5IlDWdxQpLkGdj/cafIau8nYs4q64V1cVT7zMQvZXExziodg0vrlbr86g+q4NdeJ
p1UZg6U9YnSJVVFV/Y33J5onjJbGzheJ2RdRX2oLdzXcDoJc5EGXTxPDWt88Rt4h
e+C3cPzZRKhikyhgTsm9/WpdfzvYXHIBt+d/rak9FPfbmCCzhZKTfH6HOQbaaqkh
RbbGuGcp9OlnCseqZMkhpalaLmH1YoLu6iyyqIGH17+ijG/V0liZbBFn1QHXv1Sm
ckRq2dEQ2y6gT4Bv4A19XLOnD8CUBEjXJcpP77rZWrAygXfifeY3V0sW7dNChbFe
ElRtemmw6kfsferyhUtQ+On3290U6PNAZOR5CuMO5UXKxuXTtfBwd9KL4ii0e7G8
d0S5Op9HqsHp1n5lBO1QPBqcT3byP3+Upgh7rM/aZPtL+/OnyqiLWsJA3rtNBoKh
FhqKpMiSWn8buCcVrrW+4Qga2yEJjIJoBGJv0AmX9XrtaTIqZ8syvKcOIo9nW5PE
Pat1ZoWrTkV3mWk0nGBECw3iB9eFxL0meB27ac/2pc1vmZVgpo9xIk6CLvI/jy+j
hIQrpF9sx3cSjwqjsf5iq+S+sg8U5k/KmZJ3p1VsoG5Hsukn0eIKYKao24J3K4Pi
WdPcekr8XRqCl/qwr6FOgzzwMnXFM9oQIB66QgIsBHNWZvBZdG2aF/b4OAUgMYwx
Ut8iaIyezZxGfSRBn6w9wTNzAcGoEMM3Kf90MhG06f6pPCwBG0vCN7+ewColBfjV
EPgaKRrHiT6IhBmu+oFPUB/L61vfqZwFVIBEa4nIgUBUME3Jm2oaZFIV0+CiDxrN
+6dESrrTP6d/mwnyccuCBmOXg9BTRKdP4dJy8j4wQavp0cTYZ+zLmpXN2kzGKOY/
AcNs5ep39KBmHHiTqqL8BbLfBYz6qsrzS00wZOrbC7Oxlp3MIiTstV9oDqffb5Sz
PqSDaYZRP850GwpwQZYBIq31BjV/AG5/VC8W0TX4O4DatZhiLfb3Qr6c7nfFcM15
WZ2aRPsBiM0jrncQMykUeH2/pM7GUcmyQt0gLf4ik2d5aDuAer+VPNlgKoOkG0kj
jInuD8WASOkSbSC4bdJqZBs3RVtyHEv2Xbp1febmK9T21ZHZOiWl7FsI2Ul0EcDu
1Wcnm0YkVbrh/2rn9luIJL4qivPk7qkKp20nwlqq2Y3YyT7W5PN93zCLEbLmQT9r
n9/c24ctikOK1o6IDCvkfcvX9ckJqqBu2bGO1zO0SdeN9ozX5mZevSd4f7pmswvQ
RrNgHQyUbaS8h/E/WeNq7l9ih/HIZeua5JHuJh20kEUVjfVHvSy36yTXNWrAdmWX
eiZKzHLH8zEaFUjhNTi7k54lta6dEXEpEJeIQmu3xr0yaWMluDVWJ1hovO6SCeJi
I0mjyxnWmfOTbUjaASETC69pIKUIaA2BcU8Lr5JjITuni1YQMWvRDH7XOMlpoa3A
oWM7vMfO7obRRyPQ6Wky/2phm78g4bloBwAOk3lQzEUA3DNVNBQbadXruBJwQPIC
h2E1hxgPRq/m281domEzq7tfRzNUTOHT4jgWmwJSP7XXrTs5ZRi+uuaGpbMq03s6
OZzhKVSyQf72SPqMDheKB529dDnwpqUGK9xRjy4GdWGSArJTMH9reWV5Ih66+SgI
VG9OwY2lk1QxyfuQ2H3ovOdiBbTosAmZe/GXVNwi0Xdqgg4ee7u4sRJe2eP8x756
OSLpHKkChFist+0Vny1GePXbNfEuk2ZSHaBjdF2a5PjglcNsPzssE2AVpXLBFaT/
4xgVYWqi5FI/vHIxk7jZmEHaR1d/NZgo55kRyxbJWZXUUYVsCXbhG3TuZqNernO6
RaVYvPygEYHB9QftOjBkDrDgZ9lTZQUBahpARwc1epUEvDtcDQPMlL4A/tVO9oaW
ONvkB7JII53HGh3IX37zGBaIemmXqClL9g37/gJv0p6eAZrGPmN0cvrwGd2cntLy
UosiaqvsBtUp2CC7bS3bMKgAzL8Kn3ht3ewUBbT6ICRQlUN69qizmHlgQEMKEVny
h6JsEbSgwvnHja7Dew31Been3GHFrksHY9lYkLWOeA7j59IW4tcM4mmRO84iQd25
YvNihcqPO8aXxStpn9Z1ra6RCLmCLDP9t657iUKsdhj/IjT29VQ6CltSJALwOtAr
dEoXETzVyv/X7w4A0qU6eXhS14ItkD81uylwMQihNfqiLM5haSSFANTPZ2yopsKU
cXaBJVXu3ylNICQ7jwnYj2p5SxReWhNVkfUBZo1rVxvBwdRzXJBnETrOixnfxY/m
qmkrdoFs2Nq+v/bD2izxnOjbiPpHsdgTrnwdxK3W4y0lfL5Hwt8cimVTi5VVKxZu
2koPmCpYzZP8NU0Jg/+d8zWqMsCC8cCuY74StqwkQY8DqLsr2uBmGaUA3UUqZ3Wq
9yJvHo4mho8tI4i24nPINgHmmOzpfiyXJSTt/ruytnFPlqA/vu2Hw/cG43LL+crz
43i9ATkenmznyHVR9eNgl8/Nedx1GdCPHHeHL1ZMM+W5CVQa2S0JHrA5b5tpDwRK
gUsJ35hD9e0pFvaEYe+sGp6kWCoRLr6O661unBkuhCtoGAHni1OcrgLcnu50r0X6
Xwd74g/jQ5nAGg8lY47tJ5K0A7/dphn2Q0HdNbwK+Gq0doptOtbm1iToYHeC31LZ
GK6qpQdTTVGtpb1AblKa2h74hxaHcx2jtKqsjlYGNbeLrsG7xl80+hOSGje4onmT
2EHfs4RQmoGX04w6FqYfa3b40AfsDu1QVrOQZHCDoFvnPM3Q55nBa+nlBL04dclE
fbDmoq/74+ixCcayabWkMQHyay5BSOXVvT/nBLdOGHlEWkq+jjNlHjbxuO4cIzLW
XAHRGwSd56enJMv1CHs5z0Hmi4YSwsgJbYljxTKWeUjKpSf2Wrmu4wWNkW4bHKyt
EUF6MfeOEg/d2uHJl8deEfb2+17xqnpn8sg3+ZzE4K7zb/fbpbOMU5ZQg4+5c4vX
P15D8XRQitcKEAj31eq530ZGoaRJ1sea1859we3Q9PTFLXbn8Kh4qAushfwbHYo4
556Kyf9f9iSkO6x7U9RX5JkEIi0g+dY81n4/K0+6aZSsSNxOZcnd8mjJTmztJt2a
aNsXpQ2JQx+K4eJP9dVPNOn6CbyiVnBcEHxxRcv2c53DvSyzjm/tPhqwc7iR/E6m
TrtA6VJZs68h0+lWnGdMnMYlZObzuVzkcvLQmyv5zv+m9GEh09QqV+uFQqe9xEXF
zj01hdXClnD6kJ6fzw5sHDgbAz4jjPOgAl8i3gtb5+kL3k/kZuHYk6jo5mgNlkVq
PfejorwoRIb16sW0F4BVryrmLXIePREYshbYCrfhuzgAupaDfUEaDhIAfEkAyGvI
UMXj3dJU5+v5jWW9EpxiE819RbLQ6PeNJrI6qJqiX9nPwdKkVEWSQGJbJKCPLBTn
ZLPD4F2KcciXuNM26i2qSh2Z/RVjvuoIP7s9nfT8tk3E6noyY2w8eAgQLGJ3IS/5
zttnEZDkVyMOHRNP/jShDB7eW+hpvrcsEkaZVCNsUPZ4FQpNagb1MSei7T3Q8BnE
nvXmUtLKKCYfTPK9WBTOH8PMe/d9Csi2HK2hG0wNh0AzZ1Flg6sKw9/zfQ2Lnhke
Q1NnzIhRpQg+gcPtO/hxRgcZE5vEAx+2m94Idoxj3X1o69Hzhq4ZTg6UUwIb4/SQ
`pragma protect end_protected






