

module channel_aligner_4 (
    input wire       I_clk,
    input wire       I_rst_n,
 
    input wire       I_ch0_valid,
    input wire[7:0]  I_ch0_data,
 
    input wire       I_ch1_valid,
    input wire[7:0]  I_ch1_data,
 
    input wire       I_ch2_valid,
    input wire[7:0]  I_ch2_data,
 
    input wire       I_ch3_valid,
    input wire[7:0]  I_ch3_data,
 
    output reg       O_hs_valid,
    output reg[31:0] O_hs_data
);


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
BumQyN1IdQMBtI66cn2AruI/gtuHAUnFAipPCT65jJz+1qHAXwuFLjdLvu98VrUf
sskGPu9WbQ32dyW2T2AfBdiomneufbNHmmHzOkBt7Q8c7hkeHk9Nt26+HKIna08X
qK+afLlI4EjPgEaWTAhIwZepxluhCozlneW/guThhdY=
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
VLAKPRGy4rmnyac0/NIlxOHUyEMrEq0tSRx+Yi4Gztc2+XW1YSF1oSVTzPKS2Vy7
MEL5Ua8zq7dgG7hkZPncbgHIDZKZj5tscYLHYihDDV9jREInDnmLl8g9orhRAsGL
Yakuibh3ysdDw2DToWvogOoaZcYPQQTCTJGcXoofuVVRo13Z8dgUY9snUQtHz9kQ
Rx3JoQ5lAl5QUSK8BFAz8jZuqr3ORdhnGlrEImNyT5e4iPxZUMAAx3LWlOvxmXdd
0rn0kdvWxH58cnqvAbjVU1b3VZAa3VJCLmZ0XZKuivEkoHgmkMT0DfK9IKCozR3k
gNUXTdTQ//f7R2sVpdg3GA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
iclvfu0lGhAJ9115K+0orKJNZWQpWWFCxYZY477qLRLEML0/9NKgCR/Evm98lt+r
Eodx3e1r0H+Bu99S3fgagpFk6EXNEt4lME8FzqetQQYYEbwzp5AfI389Pju5AdRf
BgcLukQ/L/MVjv3bk1WyfEEgrFY6Pqt8f6USz59tDtc=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
aPh1FdfQj+N8PM8IlMrvbO3tJjJkyL8eVr3S93FX9grIINybdGAdy0QuOVJsoUXy
FZK6AaG6QwcrLfqrzGAQ6NfrAwJUzoisalr0PD8Hy1zUDmBpepRpgUxCyMMCTry+
13Z3h6XWvUZeNWYY5esazkQiH3OoefZ4HFKYD+UtcpWBdqltY8hIKjUKXhV+Qw6M
WDgiGMyvm7SPCJDP9an2x106Hp32RpwFDmdBxwWoJE4wNsVNMPzDtpeUN7m/WZYK
nZvElZ3O7RQlcc1F+4olpc0+DMDonCkdsl1THqPPuj2oTqTgHsCxxSx4OS/a4VNH
zFoxQhZlRKfosdrZYEVDJg==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
Ul0PO1YKwRWxAazsyn5e0tnXSaF7c08IQmSIKhYesYFfhYyzniMMqqgOX+ycVMNk
YmId8CsCZ0QY3yhd75VQWhM1vz7ydTBJAPCsoGOm8zl4bJptl0uBPtohn/zZCnZA
6ETN24al7Ga5OtYrNc8qKLuDWdSmXHjQLZpLEn8yOR8=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 12544)
`pragma protect data_block
OHIxYnhvc3FZTTV4cEZzOLbaLQYzLHRU8txBn4bQkljWyNGaQiOkU8X1JcxrR6wx
ppHUld+E+/8Te40lVAhA7CPBpBnHVPT+wuVqf9GUkhF9beXpBulXRZ9N+ZHLhROU
Eg27Pxn1v3ft+V4sil1rAHeukNf/KjLWv8cZq12OR3uEwaRXjD1RPSlZsXo+lL/+
ipgl6ya209IUZ2uhH/rE3oBaaBCJ2r900RQMltCamAp00SPUKzNDW4Osdcn9ovd0
vHZKd7pdjwpfdxGVKTM2jY3rvRFWrq7CE+owdXpZBr7w2UXwuK7ghrORDdeq685x
Rb0HtCOcsad898vEKqTq+Qv3KQYiKPTdzrd6P/x5tW06OCXzsW9SItj1h6w5Gd1H
glENoqtCjSKqAXfUyh+oqUUx+fpu9XZAiLThAx9wxOT1KYZB2AJTdeS/j1qt9D97
xABB76edcTbDV9kkJJMTv+Z4Yo3ebwl6+Lke8qDM2g0FOdOR1+bAmJTQv3c7y0/K
Tg7Ff/je15Jpl6mQ4HWgCmvYzlrFAaXOatp9IkH1axDLZb6maln7Og5NrVXjLdry
o8qRCE7E7vy77QO5ORRETyK/ZufMKbI2ZqmNjENZkeHRivcyIYo0yJr/zaQVLQZT
aIqvFnCw7x/Xy+yf59EtYaR1Tgyj9rcNUrA0bRP8zusC5jZ9KrrlotQ/8h5w0Wmz
r3WHqJTKbJOutpUi9q2Q+9DRrof7g6Ma7ozjJyhuWZdcSfjZcNMkAvRCce/nuKD7
SU6e0wWJF7/yWmYughnn9uvd1mliwpTYI/1YyiAHdiMSer1AZMe5vG7X+AB1basB
TzBIM2P4Vi/M6+DSKNgyuyHQWNcv2ubng6cHb2fPSwJNQ8QnmbG+yxsQCFGItJFQ
uEnMmDfe9ht3CNTVVDkEJeCUUl4HxTqIxdzPPgaSjkn/gLKlecPC0Y5aM200bv0L
IxyCGHHW2tvMb6c9PePBqJf2kBFEWWT7jdlL6/1Rxfe614mHbxyjHxysJmSspwYy
8zvEUfvA+bWAdE0eEG8b5bxu7FLxuc2XShw1Oc/OlMR9RDMRNnechc88Tcf1M32S
OkYWyIkuSIRMvaEhFPUz/R9cZ4LBa4Zv8ISNnG4gL8BFEWZ1fgUeTaB1cBKv6yuy
UhwoTuCW5TmHxb9CSWAHLv159i36U0Of9pI/jodzEBwllHFj5Aj6n0qO3ZyUZEse
m46QG7HnvqnX/ByFbqed3sOQKk/kVbtoUDYeq1wOvCQpcsvkIycr0ZSsAHwS1FQX
9EjmlAid6CWVjeFmZ8vp12gBqJK54J6+CRrHIFhF3+5O35KQnFhirgRFSnDRgc7o
3+VthdlCZJMsL/g3SGYbiqGmk/Ugkc9YO1nq9FEBKOnrqSogg72Pd8A7T8lx9T3d
sr3MUkpGumglr+OoEjQq0ol7KlPQVHgweWGsU9WvrrEn0v7mHI/npUA7Rlo/vO00
VT/do9R1YUBtIwfJY4gfMrlpFrnaAF2KrawkxXaMYDTSa6uyIq00F7aToYnKxrq5
YD1uXc0tfK7t2JeVp8/6yPy6WxVF/uKqVmIX3cSeVLDMU691nCObzRLA05rhsdA6
p9V0pXqYsdAZM7jYRJF5p1hsavdEaX8f2+iRYpe85heaYJnrMlZi3Wng18XMtHJP
hR92IL9+HOfh9NKmloo8sS96lqN2aEXkxijucMadGUUyxvz0CvhSy/IixJCnmEbd
TxF8g8iAx55yznLJthXTT7Ssfvwuqz6Yo5MdJnzKSabrzq1x6crHXOzpEzHZ5gUH
3s63BUQRtKGr7EKHJ96Kuuzhl7VIFj9Z073eCDDeGNJieVqPjurSZ/+Gfm/ElO5D
oyJiNHmwOUlhbogZ5f4QkGS2KA6Z5N9VMdFTklaXakE3y9E2cnvL8KEkSaI2i0or
hAtOeeEHGh6E3PDKc+45TinAtViALmaWu8H5gPu5MqBieTFURsSQcEZWAlRtPuSo
xEVNp6L3Ut0dxCf9ZbwkdxB6Exy2r2WLiMkoQBDDZVAedxAdTJB0QT/cng+Cb8UF
u4KNgMKhDg0urtmJ/RPcy0x5j7wXvaB9SjCNrinD+b/YzKU0ifUcV97qOh8A66nq
/2bqIF+9aCV0KnCMIk/3NeCCsXeZzRBMw4oHvh/uy0Yzs8wA9TlkpWV0IgitNoza
sti1ODH7yhBU6qcd3ajnvJ7kg3okJjzXQls5FcQS4QIk/67UmrFEIpI69J+6keD8
ll2+wxluGqcpad04DAOypmHGaVFkw8qWYst3ChAtkBfKEiYTR8aigzooK5gCt9xh
pXoxVy7GIy87bcU+Dq67VsYIVOqPcNIokJvmjtJ5lTFfwnGdMVGdROR0Nm3gCS6a
W44GHryxPzbC/DXcAXN3LDetO0JW2M6S1t9IalXDUE2iXDBHpkwBcZyjUGtQ4/X1
bDKlFEkRZtYX7+818BfmX1d70xeSZi/MrsRJ/NBUHF7XQnuk33nYyj6IsTwyL64E
8aOWHC4FOMcccjTEOPiiYggaM9dDTqxoyci1061dvRWVIzwJKmMJLXHF+hPeFVi1
hVdNNst3x1ubojh9nk7eJKMp3rNavLfiJuvQb4CPO40d4PZqeOWigLhFingSGHKk
gjAOaeg4BNBujlOsMVj3p8tjgVzDIU1+rtTEDNsuIhQ5tmSstrQFmEuzcc7H0RZF
zP62yKMUtatWQ40pbP8NAJsYflPmlX+kk8ogdUo3ASJGaMOWDVfKxNz+vnxygs3j
kYPv9w/avT6+S1Q2Emkff5GLuyOSrn5ZjhvSdSeq0oT5/y1q1buxwsUpvXYH+Jlc
rQ3eITDhLjeCd+NHewGs0Ao2Bm0C+5m0K1XTuLqwdKtj4kvRqTjjbNp0fge0c7nF
6ffK1ohDDRfB7lExymzOksltDm2pNcJN4gh7TjHOC0LXijdBhtCBLOFdth/YP9Pw
wqOLBHyHvWPKpGxKDuxBNsnJq8UGMIRhA5ypRjzyJU78lwNJM2s5k6aEiOfKCZGv
glZlhciewV3rRSASVveIUIfAet9doIKomJvOPnW7KjO4fcU0YTDriaHk2xWkVhdX
HYjkmEypfu7MlM3RReNa3evVO41+od/SV1nwn0YYYrdroSDjMG3ONg7E/x3EEOmO
JyNIiGd/1xQQnz1H8zYZaI9S1hM8wg3K200jk4z2x4nxtHReoNj0Xe8QTNnWFFx3
od3HdW6G0wAkV+9cY38KbPNgfmxVDca8pMua6Vp1t6PwNoItgltTuBPhhM/Rpyeh
6xWBMVmvx2fre3Qka06axHg+tFCXa3F3+M5+wgI3f+zcHrNTBY4Lc6vqeFr+UXGO
U2Wni47ny7WvXNSpZ40jx/LkB5rdAzha0KJxUQajsxzAQrH5/2D0U1PncTMX1FoZ
IrAbTkD/AC3fju8ZRp8PQpB8OKgwwgXK8zp5+lpqsqdYekKHMiojFJCGGsd1kq9i
vSv/EZJyfpwrzConHYnB09fnCW+cqUeyIDmriIw1WRRSXn8pix22X7O3EQMIbP4m
OdEVKjkh8jXv7mBCLpwdfwuOWculSJ0wQqCA3tVfdvpxtH2nszca3beKlTUuyoP3
ttsbRrOuTE3PwH2+TozE4HRNrpo1MEXQLAdOrBlCtg61y0dKHJ3rcASOsq12VMja
Arw+SzlNqPxETLSPuBj73a5LAiiVVqJqp+xRNWd4IDf7TuUAc7FzdbLHtYUXJXn3
yXjYoZyC1GW4Q/Yvt0fzIt252RohtfGm2HCdtjsRuNkfP9I7YbyiJloeI3mxj1HX
AU+d3Tr54hKaIomHOVzedvLeFeeyfBZRsOaT1WBVjtPaV925YtfIzy4zI9Sv3TXH
FuZUkBoBGlbLjJt+/h9Gyl3BUSPfuYlrRFUn2flk1bonlmQxmygKkIaxAv8xwBRy
XYf8OeYB3Gvok42mPGXeSwdccvDXg8NIeYruSaiZMNz6yccmiMN5+OhUCbVPYV5Z
8FE4W4OXnWouRldqCt/C37gsQ3e3ngiCOCfQGv5LqpR0u0besKZbVoYIShcmx4iw
AUSXz2rrQzZZhfXgrOKfiWqCajUexPF3N1EcCsctAOhqoBttx35Nx+ByfQyVvGEk
/ccgmTFQi8scrcgTZZKM+sDV3xDCAEpfXRvCcrK4yk2U4sB5vsB08/s05wsdSgVZ
R9cEQDR0H3i3cMpVnDNfky5qMUATOiWyhdUKHIeJqMLxbRR0VH6mFej4hH7aQQpZ
OrD47RJQP8bfP4KD600dQE/1AZsoTIS9cryyMTlQlmf00/X6xpyCCouZL8c2bRN0
UMDNA9sHWF+5R5DzrYVc40RAAMPotcIlprKMOfw2Ki5g9CaKSMsWUo6PVHA1wOHy
4sxgRakB3xOQnTPUGgJgWT70e2LjSVS57UGPF3SaWJdLKQQq7pzDl9xwh0z+Fe+y
aAclroU3zJHdVFENwdzuTYM8/9pXvEMJJbhCx4yyG9Kc37Dn621LASsy2hwtkBA8
shqbPUNRmHqZcIKkOcM+vXk/J9fRA1umXNHZJd37us1tkndnupLoOggIpnp+lNJ2
E5yxlYBkaO/UrG7WHi6kBloXt+5OZ/xWzqicuvVRR3OjPiqa/OI3phl1eG5RBQMA
ErcY1NC9rtR46BFkYoNA/UfYEnAwmSqCyHcGkW+S9CzbAwGmrrk2zrD8dUuFL9pq
QZhGlH3UUS72mC04xnqppm89g+63DgncWQMBLphSsJkFJz6eitFvrUqaEl9LBYc0
8mqDJl7ITlz1tliOSnO/zXT8WzAiU6fCjEp2ytePSewETylj3HTn2baoH8s77LOU
cKOYXVrM03fPUSgoDlzaPH7aIDpkpxBTmLAIK5IlZSFQFg57Z28Rg1hp9jyOs6un
qjNaqh6KkmnFgzhk9YAxiTFky5mToTuc+FqKJoIKkSnJhaU/s/ABlRNfszyjgeHx
XTZIehHgJBpG2Cx22zeK8v8e1FyzLtdjnG/v5lSzEmaVrG2mp1JCFb+QVVIbJodo
hgRED5U52/aVo+wS0QUW0pgFxPQAKuqy3mCZWO3YBbytmdWZMUuEf9AjBMr9OcHo
ZgzANgLspDnIrpTsaSqXNhoD8VLpYR2A+EuJMQfCVj3TD30oo/dEP7n6ce76yfRz
/VWGTLAGmIcoOWCUXSdiXF1IByzmiUha2jQx/4Wlk8J2ArLTbJbTu0kbKHU9lg5u
k/CxsifxRiUQnATsmafzm3juNEapZI56lbCT4j3aHBFFVOLXGmBj4tuFkotd0Q65
fwABglqGaVShDnAzjmloMac58dRdW/iDJG7V6tS1YEocX9Ec7v8y2yhIJGTuMKvW
NSi+YhKEsBD7LtIJ551QUc8vDjePgM7pA+HRPnqJbfMeE0VMg97kNgHhkkoZBwGm
RAfWhJdBU33GOOodnugxnl2O/uEWdp6BuaxknUdSl5/QZJG/qirJY6b+9hpdbKDE
+ueEMtCEmgtXeaRlRL+PtcF2trR+66h2n27eOwDIBS33n0kFAglQIQ0ARxFYGr41
AyQeAjMCepkHS1MprH7SItObGz5XbmrO9Dh/I0J30XKov8gidpzLLCFnxk8hJTBT
0Pd2RBFupvtBFgPBmmrlKu6Wld4GLC94uUVbhcW+OnHsF7/k88D1+/reEQbNybyW
Xo4/tj3/ALhjXa1s1rDeRGKf/qJLYSJnZ3YYOrgystQv3LbkybvokzP7rGCUa5lC
0Qutaa6KAqKInsHyePQcm6kb1/iId4MBya6U0Mh4ZraiWG20YqNtSWABhEDDaM59
QWLB0t2aCECd//o+tqCt3efUmgO1wCSqS55LlwwwbzsTTRXwWRv+M0hJi0z9yZpH
lqMogyy9myQPDgm8mlzTrzfB3mjnyK7Bn0Ru0CigFM1hSSnwNkMsjEbL0QQiPAL/
LK8+1KxB2f+uz9pP5BBLCAvKhK00oJ77lsUY6ETAnvc5pP/e8wXlG5e6371WwXPv
nkL4Qnx4GCd8dDJXmjCF5EWiTLDO6PE33Nzzp82T/ygcXJA1NeDVggFn2Qp1zlKG
ID3Txo2UaSg5QCz74ciX16MpRD7FaOwLtMZlf0kyicMQrZw5zoNCzrNVdmJ9LPFS
h59pwT+PwlBlrC0wyiWLtQ7IOD2Xt/KWfSW8eIATAlLTYswjOiXLMoW20NMvBMip
1lMt9PMturIuLRHB/Vayl5qSbt47iC63MgbFfjBpNNSOm3CnbSYkkbPeXgSvRznR
G6P28ywd7Uy4xRG3mymq8NBW39Laj5SCT/1HFajiq54xqNKmuKZOVZza275tRiPW
7Ndwv6FzDGon4uxpYyDTyOhR5mtYrOPiUcSN0aLMEgliaNdVo2FRgraeuRg6xCEj
LwgPIPrp17/wYMZj1MUusM1QvIrL6zZEwzxzBgAKxeoht6OwCf5oZ5F/OsYbLK4u
196Prj8bcPFL+/9sGYI/cYjKdA6UADCXtynhBDR9YrGgxOVIGUhEftwbes/cJGHL
v66fgC/IO9IMXrU7GyfIrxFQZ9PWoUU4njQNk8XCsfov3es/GXfCkTXh8tD7DmT+
d9BOvalxiJraKaThQkqmGbrl+vCfYbc+Q/UrfqOaay3WqzDiJm6EEdwp6U8Tjd5K
u5T65YnHJIH5JmbKVediRvs7/WOma4DdN4MrDQ2s+ofwqDN2lGgkPC5H/Fiul8wy
YY1nqNd+PNmCd9gjjAGst5k0LAxyR8b1IkZqPMxoI71H0E4EBPUl1vcMInSAUp7+
de/DcyYrPcrVL9vpOlAqbtU4O6OIugC6Z9ohqws8jhyXeJw6YCKLORf0Hi6eoj3l
jvlCj4HCDRDNNTOicvwDCORqS/21ChXtCfpadCOIJqwlczYWF1Sh/mrnw3DlYqOI
DbhkL9veMnJEKJVHSWUvlK9ZnRTKajo/fMgJ6yFtVWChx7UG8rHLPXx1Ahbkl3K6
fWaoqkV14rPuUX2lAzhPWY1WsrSHk3IvfJXaQd6rUmJ3lJxT0SYnvoan3X/eYI4K
J05AyEtzinbNp63ba48V3Z4FVESV883Fw6/RnGxEcPJcyGfYJznoTY4VQ7IRUcFl
R8fxV8644yBlLPIQY0U33CyUgiCTj6bIxbhRZ+E0NnZPndcN6Jam/rC6eruwNvAS
fzPSlq/Gf5jRdk78LPDoCcuYT2z91hCpMpTllJAisp1p3ZluQbzMjCFDv1k4DKAk
NZePbwMuvviocx1enfdWDvB/3e1If1lPl1XSm047BmipwoK5HZ8gXy+JTLgmW77E
EqvpXWS86VJNmfsP2kRMlncMfx+SLSpE4yqR3ZhR7QePKasTL3RWysFn+hGEMIGs
3uY5ocup1TEvTh12Gfz87A+rjQAX//ryqjNdTww6n2bjN84QvEuk9XKiEiv040vM
Tx09Iyv4hK7kTyThuQ1rkIg+h1yrqyoiWCpEyqRvjpG6nPxN9gZiPsdWyk9MZJJR
cUqrHbgpoLtnTBR+7jE0wajvfZsudChwJYp2CWeqqHOwRRxfIlOR2vF03YrbYUUC
mCbDwKIWlJMzjkb8kv+nd29Vbb5wOVrUmbYo0RyNWxSqrnZk0eawAsIUH//LqpND
PvXKwIcyNpgZ/Ki/qr83GWY37h2hlEOkdB/CRa1nCycm3CgttEqgm9aLUskbEciQ
qeRMqbu2IX5/QrAAAMMVjcEV7EI4lbQdLbAUS5A5pN8R1E6uYUIDtsOcjzvf5iXu
3NiaE5DP3ZBndkiy6TKxhMzE89qRqr9DdU3ln5/xWPT4+ddbLJ54pN0SIzDWSJPl
xmv+OmBBnK1V81PX8l0QjC52/uL04bSsiggkTPMgTWaiuYTWkvXZNceCMJGPp4hj
0B2nufKJmfF1TuoI3yU6lD4SmtlMMs8uqWk4Hx9obEzV5+/w8SCAbO/l1BzC0Ra8
3DoIEq67hdczItj4gachZBVJV0DFS/cie/7OrDguS8Mv5CrvBDcZ+HcxFLCxPmCm
bgAUJOExKqsrtdNFMys/Os623nfPEMfaRy0FlWcUAfwiLNrWcxgCu9k+ZIJaGO/Z
SPthhh4czyNtIuJJEq8O3zqhQ2bwvlMGUTKMN+fhozePIjH5FbyLga4mhVldkQyL
tRL0p1tPTKKkmLQlLK0zzHwuWX/SIkjj4y6pBnGwMnPJGhzR11EYL/Aw7OgIqDLv
nua48w/Ar9bbMlKRlUIBYj7S7ipLr908bXieBhzUaVjMtc0WlHFZzkZMdQcd1Rxt
r237FuKQKlZZExSKdTPlTzh41CHtbG/K0S9/rdNWRIJ5vG3a7evJmZLetkDgDOsT
qdipYcG25lgVm2gCdqqRoUh0jnRdf0P8R7Pruhf5P05f0CL203Fqr6D6HxlxYcjK
dvUSK4XrefTXLzVLtIbIcCd1rKZlLrm7B8Wrgz+xljwYSo6tsE/66E1MzEZrHCf+
lRkXa2sb3YyyBSb/YP3MjBeNwLNNpl2paEh825QEnfAA2d0DAe5IrGO+GN+1y1yE
EWFOOR6M40ofrevaFpn1JO9P9sb99pBPPc56Z/xS2SZ+ZroyRa+a8AreIV23slDY
pkG0jwExfv35xYyt7tDTmc4vOozVkDMPz1ZEXcg8mcH7wwOJiPyViGmdn0pQlC3a
wbNoYyehSeYiZb8R6wOdKrnGB3WH7AzwKdYaFvosd03m6OX/Q4RU0A9/XxJpeb9O
5GWJ0k1HqhIsNjROx5us5R/hXozoqw3KJqP5l7R0h+Nwt2/cJCicruPZEln+/I+i
MCFGb0zt7jE1/5upItp1EA7GOs94Qjk0OkWmHywCPEC5u3YYRVxcFI2Y4Fm6OZoI
3R8nPi6HOWgziKR6gXxocuVPC9hc4+tiNhgYeib0DDRp8A6A6yBuAZgEoiYqz30e
nUm2/jYRHHj9Ns89DH4kkHOGWIIayZ/IzegLP0JUagjfJYDK6iIyi59lYL2I+21G
7F5XaTxMu/CGyM9FDChGSxbFYAlhefnAWZwHGyruDwba5qGkPtwu6JrSCkpn8jmZ
MB8oJpSe1w4TUSSvLqomMRhaxKv5Z3oHAGAM/YyXl8lcIxf1bY1eHr/em+gkZ99v
BAnhYQDYFIt1msj27ATI5kCdfoFflOzuAYeBRiLBaibZgyIgO8aVgiz3dIwEfAEX
hC0F2A7mPDQx1b8OVymu2qFf7EOCp6iS5jwShTInO1xrJMRN4etEfITyT5wS3foB
V99PzEIlwfmjsIxLO2xK091mKWKocTY7GKwzwb+jX5gXEFfafiClBrKTHNpa8B1v
j4WlM96JKuKUU3+Jug2R3s49CiuOMuZaz6OZoV+ldY7FAITLNXGx0ddpYPOM4JK7
0B/jxxgePxEMN8VW4Btv+A+ABSpVgR02K6DYmhoMs/LsRyL4u1uKV1aX2MTpNlvG
DfzWlhTumqFx5XaAjhIFX/4BGow2QvY0LMlZeZIMh/zi1PEhnpex5zrQuIHitdIX
ZrD5mMqiifYLIPlofBOEFXvWSWIgarwgSe9ar4dyeRlG03D0QdXust/6DCQxt6Ac
5xIZbAfNWAZUr7xCCYQxRFjq/bzKKwL55LcC5f2uQ4h2sNi7RLm22zQT4wsOiyf6
zp17HE2MN1pC9ed2adeCowl+4ZVhNb+pC2rEHT5wkdXYwtj8fkrfkcQDMzVUWvyF
TjJSURZKYAvaciZxOPysd+LbPjC4y07kQzVvLcyoGbzleon5GTckArzF4YRDhy3A
Y64HFgQ9MjkTb79wdXWMJKTevSewIdqZERtXz6fKtMlptZ1azCBf1AHq0G2PLwIt
8giOAEBB9IHVZFJM0vbze34c5N+EjhPNWf2GlsLV+oVfK/ByMddp6rzMm+/F1+9T
BcBVKQE5wYvFIky/7rOnXnJMFwjY2GrJMLLDXWdLfTAn5QN0AUi+ACPmcDd5e+wf
BUyk2ZrPjbmz29CBTRo6IkKdSMiFJatmxag33wQ0GWrOb4fgO539uRMtfJPZnhkI
hE/UsvA18kahFqiH7750r6Qv926RCNOayMQYMktYEQse8tPSdUFvWLm3CJyNDz2m
OOQOCXHc6FgBAV/29hXbUu31n79gwZ+VojWdUU/Ajjc+EqB4F9XcFinqxUA0A647
6R/iZOozXZNCzcpOahQUEI1FXC5JBEi7FeiGMpry+Aogd1+MWQNaJI0PNgTuwmfn
PfXYIquN2npnQ043yHd8MQ6sa6SC6q+E/fj6KAVV5ecQH73S7UjTUI+YBge2DvJ1
a/N8AQBTqWoFFEuYenX3go3SkYPe/OhMon00Fxe04c3xF5MYRj0g0MhFJy3LFzI2
2c7cHcNrXql66wbjEQFbbVPLC9b5wI5wmJ+GTGV+V+RJrgvaW8Thj2MTMCu92Rr4
xE+b90rhJwIVlklFZkyMu+28rRhNAEX5gurCl8oecjzXEE2oKQDwhVRbNIYRbE8z
dPwkjWw34/RnIT2RGPA5yKVzTDvT0HVvFoNJw4cSFTn27d2Shq2QvD5C129QzIWO
tr57qJn/57NfQGNsA2OP7Yv9XBEwGJHGLaEDUNPL0e54Y33n+Hv1p57Lg9ssbHbK
o328dfmDIpexHt4/+SdUmqAGG70EKprNYmcziEE3AtTZ8dQBEQmm1O32LYt276xR
EcP4bSek4IByTiHRps6GCXgJgFKeaqTqhd1i2xYJSWrEZ80UTjwckGmkBiCwytRF
TGHIaN4WDiMhjz4Pz3V8jKmk5E4gRs7tPIOnENvODAVZPORr+4nzN0hhwTu7883K
jr8fYF3x3gqIdo1KMS6swnyhtzFhn7FncDfiBPIwnZbQAttvQBmhdmhaCdUY64Xx
Mm+l1Dx2dHrRowWqzNkCK5+2zM57KwLxrpASc5chnujfebz7hB3ULLCUoLTHtn4/
vXqx1vDg2FQFSgHIsRzGE6C1TDylqlGf4Ok1ims7qIXkyuJXmTX6vS6Y+7U27Ltj
Ca9/rOvcrcYUak5Cd8e3CvWl/AqS9wA06P3PGCW7EFnKtpePzFBZOvaXuWYYl43t
nkh74+u8h9fVi35LB8HOrpPEHyZGa6CmAkABl3OsqifQnpNy2nvCztoC4QWKdP94
mp1At0kI2yn+UBsSixfUQoCk0Wn697QdZYNbryD8wpVbwW5hLWH4fZ1B1N8VSK10
KzGE4pLAdti1V6fQB4TB2vKBXRw3QdQHoV3ImQYOXbZCqlLxjVM+k4n/TBj0PX+k
KQB59SRNkpnIPgrgSO25sZLFZq8BDUbwkElHM9I/aUHd8k0MkXr3z15uNsZUN5i/
uhz62ahoZ/d2i4fCTNhGcpLVoH19rjKLM5t/8rjbD4sk0CS8hPtlG/DaPIeQF6AU
1W/6SAYC9JNppqu+GN8R55BsiVlIE4+6ouoo89Zfu9XHdZwQ+rSawqh7nmcEhByz
aES5PFMTPJHOoFQyMkSezPEXoasYR9L0y2H23HR1q55kY+Wr5AHQdYcQSnSomhtG
y0vpoTirN+xzJpx2wn/flupwp/l+XCSqUgwqA/Xfc0bVOF5S6ScZhBxYAOGFlW2M
V9OPQelyswuqKzBeqRYwnyYyESj2u+hWMbTEvIgkHbawEZqCeLuuMGJ68nMEIkn/
odSogQVDd3CZqBJn8QXpt3b50Hb2viCt97w+rgBSoo9B2bmlDVgxU5M/S/A12/7a
9zff9KRPRwSYA+m7E43sAO3mrru338q7Y2RKKYrVYsuzMvyaswdcm6l5+64vP0vf
f7UqSnGTpxM+O+EIRs3iICrv6EtH1sGX2iPKmAi9szFpMaFxQsjCbAcxTBlawKEy
R3sbPlW8nfr7tVCBCSWxXHzAAhakuJKx3J+vGP9YoXzwts5L6MleDQpiMq1PHlsC
Vy0U85ANHIN9WW9r9nuWd0QJcAqJBRbrFSBzQ3HPdkJbLevIo7/XrvAxHQUGrilO
OCTnhvRk6GVRwfiW8ZRvMzb6P2QO03k2eHba3j9TFNoMSOC+vK67uVpFdkgZWcdW
5ipx0K1+mUrARmL2PSGk0sr4X7ENeRA4Z8JAGC6KsU7Tf0AsWw8vuw7WmGWK6ctF
+rQi3j9PqnUY6oUprwp9fzhBG04CTuW6GHX7xfQ8/uX3EZJcF1ch97QK/FSDf/OO
vZSebdPTIjjr75d7ZhR46F8DqOa394lOqGKlRRpXPk+jubaexH0kS2JdYkD/S4UV
/hbVPcJHHPrHO4QvefRqOFPHCOnhH39GJuJVCDDUbcAtKYpcVzDBtMx6kPqyfJo2
HnX6qBhk0s2AbrR/dGKySkdMu/Zw9GWLypruf62W27JzancJmJV90UJfzSm6LMPX
PodslCSdaXMS18n85DFjQ2MMBa8V5sCHfi9bHZA4eHS2YDC++joNtULK+AZ9zpqs
Oz92eNOWc5HfYUk/0vX3rSZ8sBCDS9WkRBnotuVQ//GlXS172U6WdCm8A27ESjfI
vT7XgpBSIIBVl4fOmFJKL5fIElI+Z3WdIIoaLQG3SHjuU46ThISqiRXz2ZxjPTXc
VZ4gbqPHWdCDykmu4aiV2u8mpQDBVBNvWLGrSoht2xGgUM/pFaga7VuqIxW9f4vI
Or9lEgVqbDTSNDEpMm8UGbOd2zUBmAOkveagjFjXpAXet7cJUzqdW6s1NZMOMFrl
KeN9mqcEQR72bOHaELXuQ2iHGGwIGlfVtEexM/0AANFyVvw9EUxAzmhUGp7cIxYx
fHWXIEClLneiLH8bQqkF2ImuTHgmj10cDcG5CZupCwIQ3nYxg/8X+M/JzADoM9rG
v9OPuRr3bxFGV81CTo6yfDkImAV3crt9StVavCbN3gVUg1z0/QGhAuvXGQcDZSCX
YlWbJba2mXFQ/b9X3QZlfXXJY15DEssGWiUcPhFdAXl6DVLrqPgumAM9nntCJcSV
wCAeXw0MsQtlmvJ/LUfDI+FEhz3DJrFfRk9VeIQGkRBqYT0h3cQwI3kPUSY5W/SJ
ys9QDKPiRcGlYmdB6VrWpThC9GQSc8ixxUPEo6xCQqXEs1lRG37OCOVVfTo3fOpc
SOd1+qwGMFiAAiKJU8ouHozvAlvuR01zFzLOPB2G+VzWWeRP3DwUTHaHc1L1yssu
DdQV5wPeurzjOJEZWI234pteoWPYPt437kEA3lJ5kkS1FpCZkGGrJvP16ZC/o6gh
IId0ZWpRP3xNyfZw9OaKfEXZtCXnPYs9BWG4l+JjqAD4tLtSRZTJ9IXoR5VdPKf9
CrR0Ei53aVOyuSrMWx7Qd60xvosKwUrgRWkXue84hX+8MMH77zVLSMz05mH2blbR
h7ecyxeKRZPLURhBabfColxWOFmjxU8r4Mp+myRN67yt66gtwK7dNYQ+UWu7JF5R
k7Oc6TdCLY0/sFgKeb98A64DkMgU+6BpNt+y+mpf86fAEnqBr/0sKbcN6B7oUZwq
Oj7dHfvoY9GZy4klnlRQFPDMPbnl1656VQyJ2cBZbw5DQbyeJ8mpskScEyoIppOK
Fio8+stFx+yEXlfs+jCFY+eyuNVTxwEEB6gBCLKIkmEs0SVERMQymrJEJbtAyfa/
YNEYH3CkXPRTZv2a6BpBjSq3Y9xpidkFdk5RY9VFnxT5pYh2faw4w0pMvN7+AsWT
rRbt1JQ976WKd1TKJ/TJSyhpek/aDEu/bSJ+LSZRZVdZCXxsNdT8x733glHt5hwb
PlRMeiY1mZVG41SHsjJvi1x4ReZygmPa64Ga0S5FVwMDLvYNIj6Q6r9//rqajG0J
5/qgUkw7gphGKmb4VqvUxeoQScPvJcX90kU8tNnsLBAADQVLrSj4C1DtxxsgYnPF
IQQqJ5EJlqS2gBnQiKPSmhvFupl27AHaIIARO+s0O/cD0YepWI7r9PHNDY+BVQtH
zsL7qaQPYBvW+ku/snF6kNtenwsoSxm//n7subCDZfcaiX7YG2yzj+dlo6BV2WZv
VntUe+pPgjslsTzknVTtRlA0EOLwdP1HHXR7FbULboWkCJQNcYhoXoWw6UfnnMSN
nIEUJpR+airmtedg0kgn9NwpCIGSqC+on2zCx4L+wTbGC9UoWgH/IbKl0Vk5U+sF
7jmJNMdoM+r1d4Lsqnvj0R7BuboV1DANbdCcq6SXgk9hEEccF8fFBUyvCfJK/jxh
wtB5oWimZ8RP1iGULynuvoc59Kpg7R2tHgtNjOQRIRmTNso4jQA5+ofvjZmU7y3S
ZkCgU5TxWNWl5nXSW1MeKHDb64PX8MXGzOKw3HqXg1kDxsazUa1maoMrMnD0P2lm
PnwvrsbFgQLSBrZME+KDhmEsUbuJF4nskyFDuTqMOcNuXbHEDJi+KIe9fSClJG6Z
8/D61eoP5GusnKeutKzbNkXCeAmdF4W3SzId0gW3JSlYtHgEteOdb1REWOXonbS0
Y17qWUnY/60wQg4O2pv79ZKKblNpPXVO/pgW6354g3CgHL3ghi5G+EpNi3Qpy1UE
hrG+czhnkR/VLab6YOwN+uWA2G0q82ZKvmrGcsuJZRp7FofUJyMb9L3m0yXc7rx0
QB+zg9S4he38IqWT1+xEpq8shedwW8rz8B8KQlp27aWxsCS6ihlG7i4rzc5IB1Rt
oEkds3WMvAd+2Mzkp7yD0BTWFij4H+9lwrBPUBtTgjAUbdrdl2fCzjK8x2EZ7ySq
PK5rxwq7qJaVVyjm72thmH6aEqxnF59utFinyTXKCzF/NFiojuZmzkyOcbucJq9S
DruJvfnVhc3dniOXY/NivXvzF4PN9IpUFUK8dTWvGJYCWDGYI8x4uVAZ+xclh+PV
fuh0zZbdilnakDydM6P4AAs85wftXncMmnGDNKowzsp2cLW9fVljAopQVkSvsjES
pN7GIQTPD8ZxwG3jujPutUxFlV0HqMmV/uzXeDN4F727ToEUV6JdKxbwIwSZUEIW
e2gge/6nthIATjI0VJzUn8jqTj6cajqBmXajIxd/XXMGlh1zewGG1uuCDIrDPV2u
imtIrFdSmNED/KvSozRqB1eOgZdr6hxOhWOux4z8kP7Ge21mK4AZBHeJ9+znn4UB
sujfKRW9sDh1N1S+iebRINhMfieMEYuUXB4kXy8UlHrwgjqMFFU1Pq0ZXXSJ1mAd
YEVDZc3qQQZqpzga11id7r1XFSlRZAhQQwzL6k1od+wxyVRVPrlxvPRxugnDrY83
q4b3Gnh0NzeM4TzMXknS/UnWBaYwJH0zorHYOmn1et3amKuS0SSyeUUmWARKo9hH
HvH/BFzI+ZdmQ9N6RpLcvMqgbV8itdHqaVhD0TYc+MzaoEG/lk1kzjCPuCjlU4kd
uqAvHSMeDKkPRJp/w2ElAknaFtuays0ZXEkPIIqZ/j01c6t7Ir88+OaHMiraFGlq
Ts+ofRKDRfEKsNbHVk5UfZFhWSwdrvl01u3qUJzl1Q+Wy37hJqYDCc3JwgeeBl/C
XvLScCja6ZRaCLVBC9ZBgYJE30efJHHe1WdIkvyAxtYhpJMoxVSoi5BOW1pIptfi
kvlkXzZLRw/4aRtZBudvHWZx8otQVBP7KsfIN+9YPrjbyCY8w2c71uNTO1ywW1O4
5WN2Fx6Hq83Y78e0bmzkZ/PlqP8KGGzIfdkDOy1cArUYRHjTgI/lfO70a9LLz7CH
pjDZOwFBwVN+/+NK6lMB8sXL4s0SzWzyxHlz96P97uinbgOle0YiruZoHyGB4GTg
6Ok9t4UD6zsZd2tVAfOEcVxi1ie0Dis+E5M4nUbMlspo4/A7X+IrkD0tgdy9jSje
MbxxBUjXudAM/1tK2TCh38athIR+3CDVJL0YX5AbRG8qmfyTACuO8nv62AbeQpvt
1XO1GUq+TPvt6f5C0b10/0FlHjqrjdoT6Ns6RzLuKI5EC7la5VWeec5uZulDswCD
Btfr9JBIuZoT9s/k3lWAAbEc4KIOAisGfP9G6YH1gvSZYrAwgX3hHtkweMH5Fr0Z
BTfV87KgdWCMhHWe6X9cM20/tyV4HXEZfpPhPBWthWZe+orVz2EVRI09lvBwid0W
CDb6zW0lGJREmhV79Son951NBEjoRPmMUjD0oPBLxlggvKtw7rqoDsK86H4AH7Hk
GKOXFexbV6f48yIAs3Es9ZToh/l2KQHWRVavVzrS5YDfK88WZ0u15ZiaaD1eZhMD
sX4k7fuTtDZU32iHe5TrPEHSbLMZXHSA8vgnBZRW+4YckCUeeEMxN7LnpS+yZKZH
Wa9jABGkuoK0dc6vCACNoWlG6CTUrYnk4h9jecHmdelRgWM5Ucmx6K1cUVEugziQ
wQ6cKSfYe0Dqle7uyOLrjZv4ncGOVyZhFCfQr+DHgZOz0SLjS2hSbIdf39jQ4KF1
o1/J+gzZXRmfykOnf3o+JmEs4r2tFcUu6uVIfyjm5bM1SDPltpf1+JhOj+gurB0m
Or27C2x83F8YmtTDxa81mt8Pc2UDTOSIoxHnhpcT4GWYNUEfs7BPdBtOvVD4Z6O7
IyekVlun4aCoXssteA7ayfdX1UOJHA6BsuKnmaZKkQpeTFxubJtSJON0ZbNBKOPF
n9IzYMTYD6dEI2IZ7nvsoDKGVMOMH7qQXdCnaajmWBRNhH8OQqII9/qqNPSwhHpo
ursOicXPhpjZOYnrw95hI3GVPRPzt5K/mB8HIgbUVQJoHUBH1J2mWQF28iwD2WNk
CgNTf64HG6/ThAZ25qMdYfxlTr4ciRdJTXQqil2G/TtabvNyXZK0CPnnn+LGs83W
pbwF7gOhBol52g+i14jRXtEE+FR4YbPrCXlATGubgxW7qNFm4DkwRy6O4uX2K8CI
YnvNTxVCoZKYtl+sJ22OXRqa03xcEYE2/cBB0YqjPL7HWokTwleTryfSgIOHqwR+
fqARnb1XURuLVvEJAIOy8Q==
`pragma protect end_protected
